-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
v1SmV/1G6ywVXGF/ZSh4gMprJ7E26FkletSNIgYf7HIIe4Yj6QZRpPUs61xb+3y8hXMPcBDwFTe3
F6/NtTbcZA6VfoQRxU+hLtmwM3M3BANSyEVygMR3zTGHsTtCpQ/guD1N3tIdg16PVVmb/ThXNz5m
nCHgMCspsLDsebxw7RX8UMsEekyeEE8figL6gRMGJVnNgV5uwMwfkn7so3ns+2ZkZrSasZum8QAN
5ieFSqQAueR+SiN66WPkJhOgUqUo/Fg8UNUevSeTE2VjOSYGoFXgriJOZXzVX6Sd9ZrSUouCIvyv
HAWXCriMJItyFISNgo93A1xS+z+X2G9EbFUzug==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8560)
`protect data_block
4m3W5/fCOr6cZig+A4tO4rzwEEbNWbcec5/Fbb7LyT77Z2cSP3SO85Sz4FB0F0F60BB4gptkW0/o
SIcOaqUEMxiZYUFbO8W2jOmHxPyMsEe/zxHr07c/lNwSyNYj3dDfU/fuuVVN0LbYV35glF02xZ3m
7j5MWMb9WywSDQqMbms7NsfqxNBdhYoNeV+vquKHUXLEHWKfDQWlTS5dk++dbdydONZMhmxBeMSn
nqPiItQZ6ZEianj+Z2AFRhfK8f/yZupHf6SoHESG1V/htEZaXBP+/zYtJW5+ETZz39qGFhh9v8qU
fBPERD50zZMobwfSUFvuIiHrMLUYujSgoo5rrtTA+3jnaNhYUeu8fpQfjtgHupYw/QFfKIW3S0XN
nEPmofFKwN6Zr4F6Y9Z599oWwCzGe1Bder3PqlFJyyd3WrCmGESbrHWTsgUYYsTquIZLBBYP9/OJ
NslCshCSkGhoCeXXiOJ/wRdKMRc/FaJoALduHK1eo/Sm0gpS/tDmcO5YkYJk9fxxl7xF/TUwkAjQ
DHKqeYkKEcsSiy/V+x/mMUnHB8UiTEeP207qLvEC2ieGem5AHW3RgYaSBpkjYQsAAoVwlL92d7it
7hQORrZTPhQUM5aPFEKpahI8bNstP/Tsu19yu34gn6HOPYARSveKIf0dzkTwEb9xBhywCPf6qhl6
nIzkJ9ROkoMgPb9RAaeneWahWfAb3Tl1uqPgUkfT3x/RBoy1jn54ci0JmEuf1mG9629dzmyxhb/v
5UAR5SyX7FjWQloA29b7SkcI7hu9oC3xJFfOQcJu083gQDT8bSZ34deZDTvgM1Nl86RsShjGQGEJ
l3AtrYe0j/o5VxMGDLLihFnDAke8YtNVnqYA6YnbDbyXR+MNtxbDfAE9XcHyCNS+IhWBpUGuI6fC
LsrgvVljRVQ71UXy/9qXSupF+s6/3ZRhv/e4QM/rCAtQuIk5vDxNpBc2CJii+C8bwP+KxVt0yVFU
feCMblpcklCuM6jFB8ddU7Lq+rLP/UrSgTXzFSmuPz1SOXJKSNKZ6Oz3iVceCV15Ngm2GtqLtDrG
AqNGPRl6Ylc0/h1xHV8w1eBsknv9jC6PvnGhZBd2qTUk4Rxi+ohB/WQreVK3n9irvv/pqB7ZvO1w
YcUQd3r8qeMBcWpSZtskpgzyLAk41p5Tsx6Lc+KlYMblxKMjxz2TyIpSr3GIgigbduxIRFewGJ0r
JE6MClwKSDhO9NiqwAt2VpHMQbDRKPnCeaIPhszeT5cKZMvHvTHGhesf0MgNaU9vZ+rp4ADYTgRG
s4yPTHxj535Fes7NPVYOEKAMdta9BwYIV/8PZCmZDHWxUT0a7yUavu30qWqPzzc273OZqqSQ0qrb
WnIVuo9AXsjlTk6SpS+iYcJ1BLy0nMIAlcNVAFtvzJ3lFfd+9LihZEu0i8euJs71dmEBQeVukxiG
l24lRqRtmUQZ4ES6IeBoE2wIGBZKcJ2aM67C99rXDT2s94rHz4kXRdV9O7HaX2jpp7S8j/E1lyHK
Hs++qnDt+dmAJzZTeKiCkse0JXNQ9qpGhLoqbLZz94ADuZlOp1IQdqQJKMC46j6Zo4vHlxJFBJGV
9mAzfbHtqOXNz0KUBFpvfcGQtPOPvfnYjyTtFWeIL5UyNM/2L0ScpXngRVmBH/MVI5yo4yk9GpQj
xOKbRRVzzKeyYqEE0NSloB3IB/ONJI6eK4Iz8Zp2HHKsWNSE7vZNk1EE6uP/fuTn8w7qkY8ywJmD
SxKeA+n0joAOYhVxTvhsaRuwfQitwiACMB5B2ndef9sqxFiHCwbve6n697JCS1vnySFHtKxfstVT
eJvXHPbmgZLCHUKbgOrxYTs8tDASLanD2wSosK1FI7V1QSXoSUHsV3m8WRSg2O5H1Mfyg5XXJ8wG
zqgIU2w6XeE4Ht6POjXgKi7Haloml3kJSHYFKHf2dPmTRec0sFkblDKfzBeEwut5ZuJoSxocMu7P
M6bYhf1OU4mQ7U0kRZ0Z7xeFLAMvmtMj5jeYgRm4HaEEi7jrZ41WtsL7Y3ZjZWfHX7e81PaPn20f
xpFJlmbsFICMwDnyImjQhOd2YzlzMhGsMkT52P0ZiWwqpTQmuht5m8lSn2KlntK7iRFq4dt6jZ3N
ccgZ8KYXb95UckOc8SpdpQ+KcBslYFHAsgWvWng3cbSIT/foYIK1KfckB9V4i2PuLR1s+EogqgTc
yyg8W2Q4qGUse7+rOLS+7lFHMgRkz7eOzRR6h06TR9z/3bVcmttd+UR0ewtPBg+XOvlGD3/g1VRE
bw3aLtkYRULAWQW7wZr7ueASSNkH2mseSrlawlNCq4zqDMw9KVLKupymX4keWwK2hJMvgXMOlj28
ZsViH8XMR61STtdKwc/fiTtDqcKqqpwybA+gDTnws2/oquQMkao82m4No69M2HT0s3TYROE+HA8U
lcY7KRZe3mJOS5YIHzzTZHd6ereP0ZjnqEkDTKQEPxhDRAWrW6hvkjvBhBbUhj0/EikKJt2htZMx
uoPE2llej0Xp8ZBP3AaXXFnmjUN4xu5qa0lx7+mn2txhJRc3aROdu/bIgp+wc9Ls+7AT3tFACLc4
5d/T8aNieo+HgpmShiSys5LvLoG6wWLeCgSB9gjJFCGyQA6yHufrKRV9bf39UKFl18Y1GnBIjHs4
P41mpZqQtoqfRk2DMbqn/qXxRo6TEKPQqm5/2Hoc5FLMrSxZNCxAdHdaXkK3XF40PFfWg9PVRVL5
V2oyKy5u9qvDQzZ+DSiEFIgCQYu2Ckr7j9SZ1FHjbKV/3uI/s0ZVtECmBiSz3JjW9h3JLaR/AlVX
JGdCUI6ZxvQttFDtylgHMMryERJG4YDNu0YBHm1I93tj1JRrfFIcG53DdOzXqk7l6ioKS9OkKHEe
gl/q/EGO6A4cfbxJna2glT9vET0FPrGhUWiBawzAdkT+i4yoyWrVTfkjwXNmg61SHLMN6jZ+qwG0
JOrtdImKDObhum1JIucjMeiPw1BCTTIRC0of2HrENrDMkCSQ006aglYhBvFAZvmF44c8tMnVw2On
OHbgY4l8RarEhf9JX4vXwjtuKFzn7tQeddjqSjQEy27kDAxkuBvSiiHyBWkidaHIchVedLiFD/NR
6ToTBL9EYjyyh4XRbsIft8xZVZNIqsro9t82SG0kOkJ5V7vmL0oc7H5YR974wrrqyFd6L1KKXIQp
g0XzZ/4egd0DD/e26VS1H5JxiMmxgM6Rfl5r2SCL8gN9UQ8eKupac9T7xXhd7bG8jy+sPuasz2eu
znVYiMYkiLbe00RJEw2DvTznGJsGJSzSonT3TYKVKH79tiwqS3fKJNdsYl2b3JT7gloTwXJIE5cT
epGlSffhXWvCf8YQNIGE53dufmrenzeLKMXebx0C9wtEu0bVbZUAC3FUVWxT7gdhrXHANtnUwUuy
nvZurN4ea4c8VKcSo5P6VTnflcSLq1uFFxVr/LXgtZNANyT0o3TZaI0a92EoBhpkvnfThGS7l9dL
AnVB5sUymMnG5lFACEWxI97mxMH6ee+4QuXJdA8VuAdn0s0vVQwNdWr0+KtMrz/zaMcW+f4hSOOd
FbWe4G1eA+qWs8xB4d0N4AT25uh++L+IKSlNd9l9XBaD0btujixFrW0vGzpm6hEgxxEk3Y6Nfcv3
pxYPPv4MJZXlq6bKw5mXP2oyMhi8n7X6DvDJOIq4rWr3jGdheB+TbReAgLB+hZLAGTREipGdGO/4
U+awZ9vOoRoWS5BwEuz7Buc90faIu14tnDS9VOq0+chSpL2+6jgKA2LqP0PgewyIk0RIr9cXoBLz
lrVGSm7akmAbSUnDxhC5FTqclifw50PXwkO76SvEboh/UK2tM3sCppmmFG0jLVvwosOs1srM2X67
JMNbQcsaRLNlQfy5ppvQYRgyZAMdtsp6LXjPqqei0+qm91biaskloWwgWIJKN1wVjohnaEqRe/ak
Xu1Ul0BIosVcDTkTs0fYsDgj4MBBT6MoorASxynrIB98BGQ3gGOeuY3dojAIvcYXCfb0TKo34TGs
LhQZCG/C2ts8qGeeCX2Lte5Uk+f64ZIU4D8tSW9b3yCsLAVtSlWpUFvClZF0FgviSzlmeyku/VEM
89v8TEWs2nMIqie4Ohvr7emw871dubIoJawZpkyM1x/s6fWEXDBWVR/U06QeX5T8tV1F5iqx9t6n
MV+AdYlJgHryRchvQDXvw+RBBpzypotG2BA5Dsk+ItZX51JUz3TJtWoTK5P/Zad3SNTBnBs+mdiu
nIr18FZFMHeoiNNYNH/UkDwq80OlpEobsn1NRc6HQmNoV5jRooWMUTguNhVEBnISEkwa9K+JLNt3
AYF7dIyZDc3Ff+Knixwg/JciY02Ll4NnR9Tjnz5l3gaEXcP5RhBFkSvhk2Jvib1y3DTfwA99zxDL
nb0glH/wIlR9V3PF9BHf4QU5MqYW6HfCjcnixt2qKDci8VuCTJ03DULo0Ub31QKkH1CeU/2c5E1/
bEqMqs1DVVZypdJXJUrPWcf7ZUw0w1orKf8jPyig9fLHJYriEbrJt6pANMQXdoVvPwuIMg618gwo
fPZUrAbAFDjlJzN86Gg4IJriwZyPT/NwiE60pUHWax3ty161H7Aa6tePaLegrEqbUM+WDfBKeVm8
RQEhwMJxKYCgnJFdM939zY74eAcRA/IUlpXZNDdfhU/CLhJHT7apqKQDbjPEbKvSLawwSVAqAcch
H7DzjZTjn8NWB6TMqZRo+M/Hk4wSlWbXPGilqZkyme+I4n9HVkyLOWKjck5gB3hNcHOi24u2MKxt
zqsYSXW6zV9sMjvDW6M125IH9hHr5MpXffcC7/vkWorjecNrPwwwcDnmud1WzO3L1FaSlTkjd07L
EBe+nOaIkj3LWDKQHvPn8QSSLTqlKvJWeuqcYyajJ1VblZAJ6b7hYaBryAorVSORaFNSSBiTEVD7
xP3o97zb21Wsh7F+DnNy5c7kxukrS4yB4HeRNB49/QFX0vdoMfF+SpRZ3cm9isJfnimou/JGoLvA
Mn38yC5oxhb7JldDDbxWNOTrO555SO/GHp+x5rUOOUzTn6mmoIR04GySCLzipCg1a5Vq1X6Lz/z3
690fwQdKi/z9t3VU++nHC2oPK6ivuom8hMKZH4uemFqn3sp0TA1spaCrOj18sdu0XeGRgq9rE1ww
TjuaounNyd3Vaxhb+Eh3UN9ck1cRVmW6g5ZORy2s3XN+qXk5btP32JIPBDuiLi7n06ueC/qbsK7R
eNm5jAjgt3SG8oIjLU7dityXsjlwwDMquVb7LsH0Qdv4wT1OMhEIjl/TmogSX5qpLt/SrnDCsul+
K0Jvb09zK3ii+1W3zI4GCZe3rkZcWLYbV9UiIlIMYp770G3NYkZo+b+Mkor3KIaVwKrXgPLmQ7EF
DTuvVfbL5aAv2MnyEJn+gqitimv59PjhpHnJL2ufnB0zYDoeM85vnmkhacfudpINj4/IZVp42fvl
OjLepXocOGTLRXmJzZgMNOzZIe73etKki0JXogA6u+84N4Hpx5P7hRzN5y3zZ5HZKT5N5Cpi+6hu
T8/A34wLJfCR+eIt3iPi1lCLkEbBaulH3BJByzENho1l4VxFc/IWSsbWG4R0nSSe6w/ExTmktrk5
8emTtd7spU+sGe9bWAwLieCvM6fLjtzaC0SO0/vHTzS/smSXAT4k+pLDCaEit1OBWhKXtqRjpkgv
iWa9PHD9IxvwtaFeipYIRKGHpIiULYBxKS6Hg6SgWkyLVmIJyjz7HFaY5DfYElK4WFZc08UAQwBJ
TcKXtO598ucs92EJHOw5t3n34MBBcdoj0ol4U4hUjcdDEib1EGCqfR8sbybHejPUCD8qH0IJxCaE
UZAf/7QOM+fwbdTPL3Ibhd2qYvImz/5DZJOQ7zCQt93KtbTtZp6MNX1Tr8oCdQaJhD95Gj4EqbBc
0r4m+a1tNCbajYP3wK+Z6obshABXWt8aspxWBiUK8VItEPI3WzHPEmaTLEzNd4R99Sxrz/trF6C2
ZxDhhzAqAkVUwwxSVC1b3V7sXlB564wU86hBeKsRL31LHR/TepdwV0A9dEJM/o9aOkeeil3hn6hZ
UPqs9+8bnfwxMBJB8nOR3SzXsS8RTZBF4KOUdlN3akt5tPfO4dKhkN+SDLMdJ3EVQ8p8fEjqQBiy
5leZV9Eq6YImhOe4bRrJQHIkm3YIytV8U21p5adCkMbge7jHW2rNz8/Vh49Pgb6ovKtp+CTKb0s1
GnLjwQnqTlXqX4A3vB8gyHOoKOvt/vXzndkKazVA5V8OqthlVDMKZK2CI6CLrpWE4ZzBUd35AYh+
De4qRXpZ+wq/q0/rlSWIB+l6eZii4O+3aZzTJjAKzrTJ6j9cx2dos1fZrAannqFUGoiKv2lvrrVc
9lnXCbaEZ9kAE8l1fxU5EiAcpK5InC6/tF+wh67/WzRxbVHzy7DHKJwEZ9YT+z2Zip3khlyhM1cJ
OFZ4LeppcMMu4o9RxPpG56WjJMybqLusaRqiTsMlI86SAmE1cwffIldBBzECWL5NKO0rTpziooqd
qdKYp2Itna9vcrasbmC6cmZ2c4l3IXSsJu1iNGblNrttpcDUpl+4mPZgjD2cqMghS2/wCudwc8Os
1Qol9sxnvxcZtbx/gN4Birn3MVf6faZODiiK9nAQneH5k+f/uWrP1WABhiLIV5FO9BVd3DNQfkcx
IqTVdVH50DtfdY83TQDybrgI5qMb02youWm5jA2l92zXBOyVqhG80uHBwxRGdJc2HB4cdYDEqCX9
O34nwuuIxfdlK0SYaUS3mGzDMTVfelOVsmju7F/1NmoznCpX0wTJVSWS/mCDjZYtSpsPicAaOHuZ
bfvUZJutjkSKzb8YeXq3dyxpTzN+jRGwFS9+9t0A/hWkFNm2UMinhc4MHJ+qgnwbxqm3BjRjyoXq
K3A+prl2ZPr/c/kqS/wPQWRXbmL95ldxCMrbpmh+3+c7dGbRx3OmTpLbUQu3skp2axgtaaGR2EtT
AR9kx+LORNT0QE0yR4EhMN0Chkq8qirgk6LKnGgGbKSXBepyogBLRbfAjwjhXE7IMI/1AlNStdiq
pK7tnkpo3ANHpMIn+dKlXy48jjz8sx2NdO4Ho+jMu/+0u1DTVut8HymDsw5F4F0yZ63ji39Cb8fH
C8k3MRF4L8bLtomfkB1LmtMSEgUqrs6v+9HWMOcm1lGt2ZqVkMYwNWKYPn1Xq0Y6gut0HOY3lGly
OS2lQTWXgpm3nmVUTk2kgoP5tTBlUJ0J6FWNCmBFj8e4qvvnpzkT7WK98C4z9/6j2qMzhdJ+ijRw
AGLE+OK7vHXkziuZ2oxeeRgAn53uM/Jhqckik8m/vcjER3sYxBFNIR2K7zglWX4Ln5X70bWXI+ir
GEj4c5Vv2NpmYV2THMCXmFwOBRpOssUIbINDRMhO1nImbsuC3yftBL01901PqnTwgwj9Cb3J137x
pAdNrgRZwOOu6UsN8b+EwNMWpy23bCNhhPkZs0V7WbccEX2D1TEcuIOZ7anrpWR5WXqpz38VBMP6
ihUNUxXIcWui1KybHTdcQvjI4are26akfHr9cxE5OoChrhk8F14fVu7lrRJ36mtoGl6GcVjC/tKA
hoBqURP6qfraB4XNfO19rD5juAs99npXhE0yMb2nwKcmgnqF2LxqUuzuw9W9gaG4HsKuMwTjjZVG
ARxqALyablZowg2KZeB+bD2LEtjV8rGanO5MlOHnK8YIanUsjKkTesg7Qd8P+Jzjo0k1bOeazkM1
cBtvxyjDgqTPZ+wXbtkgoS0yiv+t1+bNIEKTfk6r/ljZ+H92z+4vIrXnUQsLv8NRaQTeLbL4R7Tr
uXYOgX7BKw8QJDBi31dC6DCWALXjijtJtkZKUypY11iKvz+jcs+htGleFTtRAygh8OEjY500JHzw
g4wMDCyoC31z/WVV8uVsZ+XhM7Q83HpdktesBFsjxB+v2cWcYP6bLdvHAfwA7UnAppEJVn87J8WQ
CzZBwaCCq7PwZw2SeVT07fFmFGQAZzkwnD9pCuvhcLqHCnH9hbM+NBS0kphc/sBGSS4hYxMzql4W
dJZqzIcuK0muT091CtIiGySc0zHPAGbmKxknYTX16paCQYmMcwQEI1nvB7ZwiZILMRYHaAeuqPiB
zuFu/WmNBaoAJ9agxIYaAJbuloVFMvrHyQ4m5MmHQu6bZ0ISy8bG5UMvnn6HWbh2dZ1doYCxPzPG
dWUUOWYTDzQ0BF1GaCfxWBSulAt0C2dY65kW/Y8c3h34QmB7RjP9cbQoY5QTusBm2qO0JFlo7cId
OJX3kZ4Abn9MgN6NoLrLBKJuIrSGVBuOwN7kvEcOB981pXmPMZIXW2F/C7uqIDcl9dNZnOVVzs8W
fUGpqclJlr5k9YIEq+PQgiGMQKxDIoSo7k2UF7HSf33cck9CveFcvvJo/r4RBZkDV7lKTIpPjtV2
pC/aR2FRg/UyIiOYwzjLlTyWcDFtIa0VFYCJ3GluMG4tKlRyevldaLPXppVnWeXZQqmMG5cW5Fil
Ca5UmJzNwOLAUgB53ppSO87MncLZRM4UQ46OUX00PfDP58F65bogd2OkBmX56fAr8PX77a7zwRK/
tA14ohrNivgKIVnsh8hUcqPgOU9TFEjk4juh+Qvat9I5VvGjjzw5VON0HyBAdLwlB3dIhTvoAfo5
BUHiXfCGbyNK6Fdzv8lfKLHvNWr+F0eBk045Xe9PdD7yYlsdWV/PlHIFuPIwg7583t582hJHenTI
cImrnrX/QD4Gu75GxohdUAnWKqz0WrBs5dm1SVy/cxCLJZJ7a+mqVGTQa5FsHN5XxbI9ISwOdOr0
bFLG67+HJSrhEQmWX/RN+8Vx7mjMcTOlBy2QdMhOEpWIMHoJCFJrGyI3MPUWqCYgxedjBIt58el7
b1oY8O2h8wpj4od7kKWRWl0J4t8ry0gRSnVYhpOZrtc3GuadNIwAkS9Xdxub0V7dWKJ8gTwStIRN
LVcsQcxmPk768/VSueK4s84P97DZN6Dep50GHQnqfQxCOIv2gUq74cjVPZR5qBGOTHRC+ikIAd/X
zmsghTLj6TX0xDNhSjxX9Qm4tIITe4jtHHDf4DY2/5B+xn7Jhi97m52gRNI1XyukNjOEXvx62tBG
y57L3IFdKfbtMEzd5dQqDgh4/QCJpJW4xdgtQnZa44Lu914smk5T7jgdb9+gWDHK0cOrIE/wkN2i
CiJbJTgW8+UOpVHJYUJRut6lhXzS3XmdZBLSwbA25wNSdcot844jycIyRsAzBIU9xQs508y4MdCE
nJeqiO3fUhCJzzh5ecuSBhVx8Se/JXg6iONe5umgR6ELbZuVCqWZjv0PjoePidSK5hNgFA3IIDDP
yThnhmHIgJ6BCSKHHnHXccJt6mVybGuReOw4Pw3PkxwwXiRCaO2jyd6zjOU3O/YcFMb5QmbTYXYI
nObs6/ZIYkCkWVLeh5Oyr1hO2ssRWFSiuNDZP0MdHYCWku9Qylb3Yd8utqHkJ9eZk8LuVJn+dywu
Fertn0TAX7wYOyM1Wi9VFne0wUUGAEjsYwwYy3rylWTblsQsuRboxT7+lXNFxgqApV0mk2dCfRfU
DEu5rv0bN98nwkfRSjnGVFk6S7pzEmKPUmk/qaPfvnikP/N96qWTLpUcXWmHftzviA0p6+8CJfLS
lGBB77sC7eHbYNqUrKaw0zqdFwS2qDKBdb8p6Gb09wqte/QP9aKJVWJPLg84lx6WYkyES+k8xVXi
4s4TJzF/O7EfTJWE0RtainahUWhWvXsW2dmmk05va1Z+yLuhDMgkGfUx9dLYlL5pphBQmTmql7o9
71QAMrEjleLig3WFp6/LfP0T8fTMolUOf8hDiHNhaHDsE9c5e2z/rcKXA0acPmS2uztkdL7D8zgS
RR554fzIwVvUDUfNjyS4iSIN5zoACf8yCHIGIelc1NPzfdM+edvTg2wRECEmTLs9hg4uzduTSzes
HR6BMHU75ARosWPo6zI25OaVqShVf6YiBEonYm849rYl/ZVnTsbOkA8XU4oSNzYe57IPYpEHrsc8
L58Fkun5PYSKd2h9BwHRnbV1gP9tol6+9uSzQkHZOMBEimdF1WbOaFpbSzCecKHFOZUoQa3MPT3+
VtrrgX112kj3L4kmfaWaId4kcXKJmqS/i+jDc3IN2TyM5xPDw8CpummHypnKE76kdESipFcnL9wY
ItjG/zGs7ZqExuhmZNMtyJiaGzBE8gfW9ehQsKBg4aPtwiuN3Qh81qyKn9uJZeoAXFW9zrYmYESp
rXs0FUb9zqCKKqmx5/kD1isL8NWZ8ZC/uMaL2uzqhT1m5IEO9XkjVMmInPqsi4W87yzBtbY72twj
oYR6WDqZyrk3qf5qMtyi77VwC/kjnZajs/JNu1YocdMEYpKXMrKPA8+yi2HsSAKEG4D92mojHiwA
V1QPviDl2rA8yLWuUuEN7IHGdGcepa4ZrFaVN8xcBvsEUHRtiSRawPZq2v96Ijs+0nXcgobD96+L
eLkCay33fZil9deIxylx2sVzv9SvQrI2t9fzL0nQsAupDnUHM/Ta1G01pS3wGCqeH8C/GMytS86d
ADF67R9pkQKNTcgk9lo7YO+lkkjWMzwKFn9IiM4IjvGV/ULKWyH++cNZoE2QRn55l9ZPGkUcp7Fc
89HfitL3u9vZ1R2bYN0bY4Jko1p0PfZCuxLR7DgdQ0IFslI2ronNSCghjzDTOwLheEm5VRc+pgNn
0pOBevgqRm6hEi32P8KSrjqnqnbDTEPKOozEuV5mbR3kKTyO+lUVIvEUOlOhHfRqxmaZG5RPOHoo
6rcKyrumYcWMqXM6KwN+qsgd0B8m75e2hMU07k8gdFO8tYyy1A3i5KYKr01jMlPefjiAuJFLjc1t
UIMe88n8oomn/+gcalvb1mGFzENIA6O0+R4e1oQhpnjomoPZNwyQUqHsrxmk0IvSZf2Oj1oQcjsD
ELhCBUbGUkPeK3/TmvoMHPqh3K3HV9WnPTuQGcOBBxXe8c7KV9t9Eu1eMjSz7HoLGlK9cFc7ZNmC
C23hvZCP6Yju2XDWYVB55+nAlcgzno73FxHzhJntTuWUQXQpbbuGchp1lyXsEesA4BFmB1uSDR2l
HKmT+viSLAOQmkL8/wqnehue0F4aRAe4A0s2zguc3a8Zl7N4W6xr5GH9rkQ3xAayEvR1m5rmVTpJ
avgA+gi3iNk5fNy+RqErCzG0JLPEuwB8YCdyPKanIj6fR1WcxH0wib+3NG2CS3dPc5upOkvq92qt
UbIkgWmZRldH9EmN9B4aiWGR/XW9esvFzqVIEbZf/tMi1psfgNBGnn/ap3PW4BC6g763zFRGFxLd
OQxBtijcjEsSWhcSETyq3Ty9z0NYDx6OoOllJYtc+hx1erAoWuxK0KH92+/2VOrFOYjWBavWHv+d
nGG7dwyxExUSzA==
`protect end_protected
