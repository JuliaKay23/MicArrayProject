��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK���mkݛq0ٱr�Z�8:Uq}�s��đl+������G�7�]4z/�A��cf� �M�X�I�7T'R�(>�I
�K �udK��$�s/lW�_B��tI�u�9�ZYY���׿[��B3�B�/ n�z
_��kH��	|�6±Z��ɰV�e0�jMOHE�̨�F�l��m>�gga�� ��4�8^G=��6U�2{)~s*/k}�ӳM��M5)�~a��?T��_��aЀU�;�#f	���F.��nl��wN��:��_\5✔t=�E���n�T�?0����o8�PĄ� ��m���������;�TA
֯�0f���@`�RN=:�^����?S�~�1�tl�	b�Y&i ���IO����%k�+�x��qcMD$N;[[�\�d��y��
Xwԫ�P*T�$��R��*��H.Ѻ�Sm����(�^�y9�j���� �����8Rq#.Ee�!s��������F��s���۠�GC(��-���g	f:����Н:jL���#iP��-�D�(��@L�<���TD����^�3�VDY��wGdx��Ρ-��"q��V&�[�j[����k��:/-q�5��n��w5q�<�)�AŪ�!/��y���� =��~�\x�?ݛ������C�62ʦ�����ْ�x�kߜ�	����}4���A�xR�NR7!�>�m��0O��E�[�Q��s\!�S��/2J�m��G��nǼP��\��ެ����f�Eu� vN��g���P��,��9�67�K>/�u5b^@ '2������P���p�P�e�g���������zM�Y����F8x�=�FM��CB�;<� �����Ky�����Ӏ	�ʦ�0:�"�ɂ7��N5��!�5S���3���ydEl|0`��.إ�ї�[�ʪM�қ�E��t->��H���P!��&>���b�/�I�"��"�`}�t�e/�{[���FɆ��ץ��A�sV�>���n��kQjW�}PqY_D(O���p�f�gx��G�T�q��5�FF��A�zC��	�CNl���å1������w@*F�X�28��Ref�����^��	�l1F˦�~ϗ�3ְ$ra����T�fo��>l̒/H�&��)א:�7�����ɡ���� ����8�m�A鰹B��$��E����z���p)C�����k9�;��~9a	O���+S�2v�%L�y8"��C-iL��w̜	S\�O:�R\�OZ��R$��MK�=�1C�{.$�3�1#Ŝ!m�����+d��Y`,(�"���9H��X��Y���gj��3��a�>w��_��r2%�p�O�X���F�x��M��6yǢ�q��|�P��m�A�/"(s�u�1+�1hC�u5R�S�^p=Om�}R�a���~y����J�
��=�!�݃��ޢca�̧�`��E`�]�B�
�6��K���Rm�'
�m�+��z�Q������s������g�4�:��2��=��� _W����oLs~@g�8_�R�pIBY����R���wW#��?�.͌d)a�X�X{+���r�.6;�Rv���"�����4�'��3�����I�#��B���W㧬qsk�+���4���U�1�y���#����3��E���� =�k~cI������׈7�w���X��(�<�\&نM��PO ��s���g���Vp��ɀ�������~*��b�J�(S�?fp�2��M��!��>a�U,/��r0iI8^Z��95k��!��v�����֝+Ͻ�Ķ�BW�?zsȂ�
�^�9��0��|�8W2d_�QI+���D����>���/�������w6�h����/>R�/��"@)���[�S��5z ��۔�T��V���o�������y<�B�r����몌V�n~&-B4��+&�hз˸ހ��~�V&
ۨb2���e��Y'�/�c�wX�z�IU\؞��k��c���n�+z�<^�)l~���/���&�x��tn����R��9��!80:���z���L��g�Oo>b~�p�{X����^9G<c�m���yn"�Q��yN�u.��cҨ7����Xh��)�~�w��[ͻ^�W�⣡Q�n[���+����Fp����U�Ǉ���D�K�:*�"%���a�	��9���X\d �Ƶ@�F���Q9[��/��sj⢖�.�M���ɇ}�����������f��`�锔������mD座�O f�"Q�>V��/������[��=N��J��^�%L'��ޱ�2Ȼ�cj��x��`���\4B!w���s�!c��H�vh�YzJ����<#��M����m��9PR3ʡ��-X�\-��t|��7?��bC�jw2�����5��z�i� P�o�.n<���f��[��1�d�u��{���8&�zgX�G����Zg��l_߈.�ȿ�ْX>��8�	d�i�.8��̷� G�d>՚mI�yճ�/��#E�.�� S3������:_��Rj�8x��k^��e9��\/θ)����J,��.�ڷ Y�9�wH�Ȥ�v���|Z�1�k��डR�əᤇ'�1�-sO%)V�o~ݟ�d��1o,Y�~��XJ��U�D�Y�6eǂz�g��:��q�z2@(�F����䟔�%�K)��4���5�	�����ٟp��V���F�j��8`m�"�~�Ȧ�E��#Mz�;�SA&��q>�4��~�=7�Q��kyyV����ɖ�A�z�SH�