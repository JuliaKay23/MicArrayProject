// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
RbodqV+U89xuFUDqYcAZAahAB5YZSDkDyOCGTWoLy63+F4vyWW7dvdSchANVDDypl0NSJxqTiDvs
4Dmvi1xFLob47UyGvNDBD6dkTVVnyI3BKU1c5uEWeW5lMR/21rVLrGxrbHKTZqHIZJHeOicChmru
RonAZPvav4als06r4lCMsoS+lRIrM47PYACOk6IaMJ3UWfzDh3NziKUg8PBIpY3FnaZi6Q9GnDaU
Uz13PRVGljxHH5oXIY6askZjq0Ko1FQ9IG3kZkqfsebRbvtFfP4WqleSY/RcQRae7DGrnwxIFzjR
Iy2EZrYcioVc0HX53u93jY4e8v8Ah2wsCPLzgQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24432)
kylRCuC66lVtZB7/y8Bj3WJp2BjgowoZgS6+CdIEmid+aPDfSAFAEz7vhyTxxx3B+PcWpjO/CxJp
kWLCrL9kPF0wb06MZPJfnVvzGnPe8Ev3GNDnw31Vqmoq1HXVmxkO3dAgYwlMWszjXtJKjNnxXvRq
8LNGqiWwDFafHVPbl2Dd7lD+x42iDSMw3CXYuu1IVR1k2CqJ1+eXpIaDLHKZZh6RzwgiMfj+OSz5
P5rUpayRYx6SWrVsFBCqR/ZlcRQBR8E6gKyKGLBaC3AlCe0+eDVQ1Z3rpqlZExvIX9G2OPu4euaI
llQZ3abwfLQN5axgIC83wyvK68GM/lPdy9XkgWkxiNVimlQLsVe/x5fVphs41BBnIn44fazqZLl1
9igmx9/lU27swFee+BUojWVuNrcyH1gbZzQxgJIOEj1FU7YzSJFYcrYZ5ejX/4bWTCmQ7DEs8pSB
hyX8Gr4ZF/KwJCuHjA4a7ShyUHx4aCQSx2htm1i1g3UXc+n3DFDYwgKLXF6ZPj1Bd9qf0Gq5+Yys
k9tlBjy7lrtcV2hEwdkxd2+PlXelAykpdMN7lS6jLCJMn6L3ME5Au5Mm84Unu9lDKk3AAkCluGzx
mfarXCW7bVvNxQf6jFUJ9g/jka1h4xqQU5gjQ/7wDKamDT9Mn3IfzDAifCmwQJVCWle+N9T5H0o4
7mo4lRDs3KFAgAgBsqMiHkPhp4T5IDANgxyr6iP2ef/P8S5CCA3trAzHBmqW6UO0GoEArY/DQUBW
/SssQMVExIkJsiAvUWY9EbLM3ara+/JsFKKn+zIQtG/cgStBWETPVafgairCzjIOgSIXBnp/MQIM
D42Q2wULWtqNAQpUZOdfLc9ECQ0vL7bukcSYqNlfU0SgaQoiyRDG/8DcXCCEdu6ZVi+t3g5iFutn
5LuzR46Ir3+EWAZKwwaDx+LQ1roHyakRIUK2735x+NyOyTekmVGRfeEtSvQNJmlF4xjzdwMJg8E7
2j7CeDn10pRC/fx2PVNawDzu9y/cH4ncaZcLWxRnRHP+Rgw5NpT5l+Y3ciipdXWznUZGy++WpbQm
X2MWBIaZqlWgEwqTy8TTjiluwUDzlrhltUm1uhkFT7jm0TtqDvmLnDgCWww5QcV9JmaPG51WYvfy
/BJpsP9htfRLVyCK4e2PuNnTacSxF52ZJPEsZRkZ1rUuI84j4v9cWJxmUMH9PBezWNbq2098lUWW
ChASwsskuLV7r18w8ytyjCAx4KliaIBk1P7Z1aljPZmzBc4bewLFSiURsh4KMgVwDlbuiDtmP4xw
8fLiWwvFuYYH4/66ao2uDof1/JapOufmLyax1EbdpoSxUEeMMxjZbqDpog/RtEn643scZyTwT3Kk
Vrtj5evljZqwxuXTj4L3naqkFTddGgbrQsmfAu4EzkT9djz6tTPZQTT4S52RuybYeAjuDANnNdlK
lB4CVRhugqL/I6H4brNxEI50VRrYYlvkMXikAXTN4roxT+hB9UZASYVuL9+On60jZOY4hj3mTnDy
/LkmCvOFgTJIrifHt/2/tTwCPJrEKDT+TJ0wmJXOejqC1d7bJvCcRnsPQzHO+R5+Z5uGz+SWhEMI
uvM8Ykb7+QpKRZ6MSZyMzhpqfd9YIpqhZBgu4vWH87oRK/zVpDrrl40RxPw2yE+/ERwa4TuhAmhh
Bu4fA2SvytptgTELG5qAb4+X+xh+jP3PrzKB2Pw9OIQ6HDaic3plRrlkqvM70Cq6cAdPotXXidcx
dlPsP/5sTbU11RnNA9r8rGaivbetpdP0fm126V4JYO6sQ0FnAh5exKfR5awqHL3XdNhOs+8Q3R9N
T53j3dyvDqxTNBHXvqJAbPXIXeIP8WSmaSQQWj4ZGO349YRHpd3Kip9nrjFpFKQLfN1ZU/6aSyuh
ciU0JSlKR+cE5BOvhrXcJBzDbAbQtb4f6ob/v0nQKgu3wlsUMkWFLixEVyVvpQhD0cL26O3TJAXa
KuS328oZYZiMxu9UdCZiQ8byqnY+POCSvtFEP2nUUyls3HmInHADjUjZ1PHWelewvP2STa/O7v6+
lGi7Z/Wxgy64itAauiOcQGPWonG2LH0CtDJ4/RR15dEs7QrThIq7g/QEz0HOiOT9ALCfgk0APuYp
KP2lLdAtnpGCh3e2IiZp4WZGIWhQeaUl7Once7e2ciUVvfwGIKdhvPE6bq+8Sk08zFU3Wwrs5YVX
OGxFobMzFB8Xg9cLToDvF3Fa7hZdtgeBuVO5hOPlmS0Id5u2wQlt0bKiIiqc6CQo/mwQMLZRJ5FS
Sx+rs/6148oMlJdcYn2UbiHRIs6fKBf1pgyOsRJ14ZAqfrya1sD4Q4bkHa1mAsk/UPfWtV2BE5V0
pWftrxH/QtWRxca4HBuMX96/367tvM9nFk/3zZdIzvV/mHNEjNQxhMYTqWDfkLvB0uKY6Mjq1BtC
O4DFiI05yXZSUkJncf4twvkQTSPHVouO/lHRcGx+cgQU14a5IN6ObIBAn94ixpIUAmpbfk975H0L
bGNfnGCFc/B2RNP0e8sqhXBuAmpMw7l+mL1S887LdezqTl1rhAc9MSoKqwPrNAkrYo9PQ5q/gPuj
0MFzVvCp4Sk+ls3CpwqEUHXKLMo1pNXChbJNio280DqhShG9wc0ZDvpT+s8drZUQqFtJGCtlb/rW
1CUkJLvnQijMBKzznXy9k9GE8/QjjQsMY3tdYtTtyd/ryPh6VV+aTsx/4HrV2+PW6in8BRK6jbeo
17TWqZRTyltYqeDsklC3WXmO/f2WyK8CR5c9ZLiaH4xLl5jq9fINY5SWsP0cUiuXMORMPRWpGM5W
kx4rM6H6l+mYegyblsYTT/lT+4ZvRlJ0FTMxPBGXxsq/aW3LGHJ9wvmE5NpJ31tMksAj61Yi+9sp
g0GwllF1ch3bpodseIlaikTjUm6BQxLd+xMcqEkErZZu/KwBXagyVULGAkFohaZS9W64T2qH3HPL
JDJkpebKRcANz24jihqLrHy2z0dftqEHL4GrOijV4W6zt0ArG8dxgOYTcbb1K/5RodM4gl8W4k0V
3waLz/Fy4lyUBCBRDgPo4mT3R34c45pNmr1GlbwfgUoYD2Ha6jQYdFmML9gTQv0sH/rHCfewal44
0a+TX/D6z6xpmd32gPQHNc3tBUZs6HQLf5ZW+riFWyuOJhdPGxMzSZtjCNtJaTLTdnIJuWeP8BET
lwwNlFpwK+KuGO0/TplOTV0PZr6ulSTVTrQQD3vihEZsVWXv7jq7PQW/Z2twY1VT9xzlP0WjKLIF
lF3xUN+NxsWKXqEn4QpArqpjYw2oX9/YHxIpx1oT5iwixB5ao5D179hH5QNW++TZQ06zXPEzcSFC
6//lTdNoKb3oadqGViHGYa+o1GY3Ly3BOuqnC1hGGYSWL3SIlpblAUf8cSpjmfFT/un32zqmCeyC
yFlwWG4vgsjTNEE/5ftCY3QX0BtKcmWe/Ocgy+lfeqxaaKRDWTeB8HFaKejuuJahxdzor308bZeM
96pQu07TX8bJl1N7bClCjRw7Zu02Zx5At4bk7hkGQreHqBDODb9kLrbG8QneSi5/SSZF3QlUFyoj
vmyW545ik4EPDnb0jMSki88fdPp94e/b0XnfLsHn53T2rUYR/KHYBIrbZVL/t9Sm/71byICfHQiE
Cos3dSkcAtayxuchu26twExvYuv54D1uzN3k8O9Z3OdH8HKMdh12BPEX1tiizZYh/8LurxptHvqB
KjP3OOM+ZddlC+wNLlJ2tjH4QO/lRP4tV0W8fnfCmb2y5uz5hU4jRifMdTWkNKJcIHKQLpq/DP7b
p4/tUXsC3/Nciz1uBZwoD1uNvM/D/pFkItfw1AtlsYqdLJe9l0H3KdZ0wvpOmW4zPkQnAp9QVqI4
hC9IvckygRS6VXDHPCa4NeLvoDJIykEU3/iirajAFj0CSibWPI0vdo/gC7dWMOtQLfLwyaXvhRUD
nAddU5cZwNbcSxBf/NFyn3odIySLOCHXTeE+aDVN+apGI0TR45sO3jTonuo4QrrOu/nkdYNUcQ1H
+6IHRLEK11bEF4a/CZSjob0cnuvDW5BppJKu0uCCUDGNHJ/J8fGd+8YH+cEUktG02cLvWHaHlbgq
6F3nv8siRhy+7t/xaT32zkNjzsImlOOfQOxEu+zAgG5uLmQj6Beew5vxtZ+scdjQ6UcXfsP6qIBH
cQC1MUYi4ZpzHo5fLsegjrllnpcjCtJU19jBbasd9fUmKc360D+g2kJNvEAa1LJiIr+FnaqIJCA5
Ns2zk9UKlQ2Z5NCLf0jDb2BOW9GBe1y8RIMn9bz+szIPZ3CzXa41V57R42uzazdBgrZcmCrj2u93
JRPVuc2cYmPDcz4gWGfvjFX4RthZpD6QfFEW35poEAtC0mxyaJhhS+O4/gHEYJy/afJLnlpIIzuy
y3Dd9lUrBSN78tDUjcqhQqyfZBrWVE2hGdLO9Y1F9c1h0U71nBsc/O1E0w3nSeEll0eHHtTGp+qT
qIGuDN9cjyXClBPebDJMGkLo1LOViVjswXDZc4N5zJXQGkjxi93WrPztqj1o3P7zfnBgu8OJZ1n2
d2eflerBJU1yD7hKmqMi3aT1zXGx/dn7Rg0Xdem6a0EFspKmT+RC/oPewWRoPN/rWJ8S9JzPAmA3
fi8VDqHAUU03o3eLOceLMWICsNZZM/enthHeAxrmOS51Fr12KRa0EfYW8r6rJajQTa8Qts3aAtTF
a8Mylfbl8DeIh/cZaTCz/3Ki43pr2QPVARPWy2KD9ZyeNlb6qWhjCDZ9EnhMtzEfifHMdnkub+u/
0kJm81NDVdkLBZ/vUeQjyvwG9o7NPToqNiRLI4NP6zv3RELCAUVf80m9S3KB0MXAzUciDRj22ZuS
dHPiT0tZYEiHsiJbJ6HK+Ze5J/jpKJA1YlE9Lv+C5EuTQSBBbBE39BcUnfVusIT+RAWAK6O94lNK
3u6jK80vU8G0Kkkkp3d4J939mOQwFkav/rZnqS3irNVROP3iLRniaAAXKF6b4YSJYTGStUGZGe1p
09w5f0zxLchQbsG3uNLP+xXeij9eoIQafcOZ6gR0atEofxjh3OKaHHzoUbhrgu99qaBmsrUeuz3j
HSzQUMhcgIobHHpTxPIH/qecpQnlqt7mkKMuCTIs0p0VPskK3rH+psP2/ShCAbJGe6Damx3yUZ+7
6SENpuNPAhVrDT+FZnxRPheXs+5jh0bdjhJoMGMABBiTD0KNb7LhKy2zrf4IL0R9RRjG1qeuG+yO
vBjqhJA7Cr0NJX2qJ6zDW+T8WMEEbUEf7uSs+MmnWWXEtRlkBau27KGPCF10+Ye4D5dBKQRclIQK
EtncTf/1K1Q/GbbcI3HVoD2DVHDw+aWlLRlH3osqJhpfzbP2f93exm+9rVk6MdBcpZBZ02Q4SPej
Jl2t38Jy2KsjMpd+b2eUt/76bSHEK3k0cQmkKt7lgIKgqzlYC5bK+14vPCVhM2oOjDMhIqVDAquk
lZYLli3tOb2VNKb/9juk5YongibW1qCPPMlgY4d1XEuAFFWC2PpmIwpQgR2IqD9fsKTJw+Huymqg
KCZ/z0zfH8FjaY52G3SRC5keBFfTFgjuCEHJTwkeayLt/xOPGZ9AtNI7ArLlXqQ5nuUGUiXyTXMw
1BM0RT6Nd6fA/NvjH2ahHHRfyTN8BUH7CDTirrOW+qhEhSRJyJOFlnTbWTmZV1xybFtXsUUbQ2hq
6N1EUukacIZKlDpAKBuqrz0qfCqMsIDdbKTK9MJ9uGCStciBluzY9IkOpnQY4nGfRoR5v6cc4etr
viUOz4TifBqqlVo6UovEr6CN/QHw/MWnHNiAmSUaH4VPC37SFpQFXwGPjoy4h9WkMRjbExj/28lG
U0jjK5uB+ccfsBNhwGXT9qiu17QBE/kn9uEk3y0vl+sZwON9rVcmtLLPX7hGyESvVmIhHwLXzpHt
8etDMK2AOqLxGVZODKnCS1bdjOyc9J4ucNFkgAZD7qOMYsHxWZbVaexRfwgCzr1CH+Yjy5Iz9bFq
urLve3GWaRgGO+EI6uryrgoV01lDARbRH3VP6kptW7a+Bi5RkfQkrsM06iQrbu0grMSjPAjO5i1f
Is6Di+lyIABCWfzMG6B8aoO1dVmaXpZDBlynHms5OA3r9itZYWbTa1AwWlt4V34nsr8UqVLa61VT
KN2ljV93ZsIcDVxbQvIjZFePJOz3X3CjLddh56PYsJwryJADEsJ1XFQY2ZIve1Rg+s7h/odHxxN3
v7ZQb495NIKKOL+ep0wbD5ODfTkVVlJhnuKQDpFAlwDLsviijATs5k3rF40PrPfGaIX1LPS61i4a
0iObtau7pyNmKN/tcmhOTESQdZ8QpKfiQLzxcJq/kYhtSCYkXq0Rlo4zcw8p3QugZUUHVfI/c4Kb
h0E2BMtEgyWKe8J78NlA8OpMmlva2FWwUTqrrNXQYAOQAcaIn0qcAR7VS5/A8A/FqdQcuWfE8kSr
BriQAcL5y1pK+4lqBGRf9lRbdz/J/X4n7FmBM9XeKfZEYloxyenLHGqldShL/D1kr9GWg3oWCc9p
Qdnr44WD15HjE3kEpQEwkuppEeEs4jBgKuC6P+aYPkODXtUk9+h+hfiyZkho8an+PEesHI6kkbtR
KjlmSZDcQ+yIy7Yr0l8L1k9MDE1H/SUTxZf+evGmmHDuAtnPRoJ8vLzebwaVHWVzIynwe5+cPzFR
zAxVHJgUmRuJOYg/ylqGQZZ6huugOEgTj8RgCfXDJuyllbBL2orgdf/Cr0CuwS1gPNowxmyQn2u6
q9Iin0xPMaC3ZSWBRsWbSeNHS00AFGL9nWDLvnbv9myygjqF+bTFKMdWiI8WefqZCfPusMQFZRsh
VVfD7bBB7IRmMReFxdsY6rB0OqQqQOjlFkog8Ss2mKpESBW3AvkRKgYZHeDwLSeCaR3koZ1Tot2j
jES/oqlpryiQAYA88hNczb7wLEE3eyTZyA2w7Fv2xLYcuTdgt5BGANJQ966EUFHBfAQMFkxLtwA5
y0tJROwCH3emaaQYPR8jwLeKJsuykn3HD5i+4hLlhxc9t+7QnpdXSItQ2eF7wqyM1T8p/2+PaRY4
2YqK3yquDbF7INjJASt/i2Rr24H7KPAlGrVrAgr9RvTbcs0QVzfi6XwfqfIdxWQ9vL9ftShthwdY
9hrpCEYX6AUSe9cMxHS4mB7BBqqrrZz9GAur6efScSFTj7rLDEPVON2A8DSauH/xukhAVTKIaHFK
WLaRqXL70/9VcCQxefp1i7zI+6DYubslEut7YDN+AwMja60vv014mcEQdrOfx5Z/WLDq89fRYEBP
goVikB1r2F4z7q3k5PKCGLti1/2ePTCFZRboX9RZx2aBG23AC/qcz/9K7BAsRUFgKSY0GhQ1INo9
2K4ieg+C4tolXKWv/t5VZd4ACHrVkZYMCzuzb4fZeyGMh/BKWXKDn1cNz1XPSCOxkhDRXMlJezxv
w68VWu7z1Z+lESvgN2XZeX3tsFJsScmHAj1QA3cggVUFd5C9rL4nMSfcU1ZBEtbo/ISyAVlK2o3f
npN1FgG9WnPBmOqC4T86RpNSciIciOsZJyZKzFLoZF3EXfCOz4zDZaWpX8ekoHjfr60fpThhxuWX
kAYkie3cDQ2Q6zos+mzkgfuPmxDJz1zwOKWHentUUD9aOko08vJc2RCmERZhzSYpBnZgppkmxE6b
VLKeawR0U+fWL1kGowayY3BxsYH8UV5cMsdy2+Wn56BsOAsOYFfXrRBtYp9tHDB+dsobq7oqo6p8
TMgmW29gjHsPg/ClMrJwXWru6Ua3eTwOXOSrQLmhQm8NnWttAXBLdHn8LZEbEu+Id668PpwKQDpC
hlVfsZMd7H8stGtnCBsAp4qRdkQ/wg9FDbOXr8WjwxQano5AID1pwL7IdIDdCR1NsyIMyaEBYW3H
BJo7pb3INWiOOmwCD1qp9GqAZni0zXsBJxgzPqtr3k4yyV6tMcptzHzynAL52fQImretNCcH02Bi
2UWeRLkJgk5DceSXw/QRqDGIE46Hw+TEWelwm+WGTivVH7w2KFMS+6peE+hP6NlGA6tMeRYbQR2F
54B3aOOlCQPYs9RQxx52zSU++r5b2IDHu6eFhbxUp79vYpdQfoFutlpcM+1N7QnYPCcAb9F5nVLE
65bZiviCKQ0Urxf74LWwcVK9Q5Lfkgj50B5Yr2HERogy8C8QnlufwLWM2lYOpe2iYkECNOO0/wJp
O5k3eToXnxSvBfaYkyHY5m0Awy07z3/GuDdwr/cjO59gQj2Rk2N1uczMQg6HjaW9SPapbwPAdsrx
PP6kk75i8gyQpS874eHIEnhafHliwbmXppXkxRBSkMJsO9ucmI4OiPfofmM/s4Y/dkAKdL+JYRFh
EAvp3QAGsn633ETZ7STDxNCwpELdX+4heB3pVqjaoKQoNpqm7CJdZtg6qEYZDdmtJmXG7tyk2XUw
0nw795+5It+zD7fFs6pvwBsZeHrGHAa425u1Q4fGgaF+8iyVpi/unmboY/G1H5TWJ3zXXEwQCgWh
A/SXEhrlt3srhtWr3TbctggJPuCU8KeabeJI3P3IJ33f9+U7pk7i4WfGuCnYlI/QbF2DfzgqobRZ
MdKnhFiQk2MTmAxPtzZOJtSBEoZy8g7veATjZZzF4zgBBEi+ykAI2Gyr+bF49YKgzMTGwvkkewVw
DMFPBSoMwMs/Lb0plSdNbaP0QyqeFyss3vbFLDQoJDNo6s3wAFX2YpXYZh14NZbjQQ7C0YR7aLl9
eeESV/9tO2ctQ3e3oEZdjF3FcsB7DHmFy5cWRaBP5UwbwJRp3nEzGk/7jqECNMNIvE2qYL4R/9Ux
ii/7zr4CGU1PBGxNyYaXueQObgsT3jYWuKRDRwB5uM03bxQ9TJnodMp8fh33YDW7PzZzcLu0O/YM
qeTXLPvIQH+/wSuD95XPU8K1dyzFuJj279Lx2A1YNZ+ecymqOJmm6z5ui9vXVb8/EF8ri0dw0XMl
dYwYNgYIkqe85hfd5lwnVqHnuZnt1wjDZVsJqZ2R1chywO+nVh06pi162of0xA20cDUBJWGBzcxe
qkLumN9AVmTRZAjD1qc+rmX+zl5/3XW7jFbuLIlzvsanO8cTEMeyqCaivqNIr+dh5vPPTMfxYt13
/FtWe+anPsWizZUskb868JVujwC7iJVVrC5ae7esb2WWp1S0DGQVOscgGZAITZpsnxU6H3MOg6BU
AlHTmbeMJWAds2NaTdwi7pcxyL73oLfRZcx94d/LAHyITt66FapCW2hKiE23dAqCNgZrAb6IUAaM
uQGU5eKe1B2SY8QZJgEzUhbWAaN1pFObndWE6wkTPZbTjmWW9dwNEHmmMhwWXuHF82TqXePjtTDN
xtr3Gmtq1HkEun1vYKb//Zg2sujrje1RZmfgf79G5QxqtDjCMxmp6N3awu57A7RD9cOwLb1ULD/5
PAjmNV62kaC1xJO9vLCQpC9xia/iYTJMP61UfFs/e9J7uROW3fD0BnX9+9qJubnRfBz2Saf9xb/a
h+quDXblp6ppo7liUB9bM2SoS5hqJceapup5nh1g4IQhxkhUcowV5xaGJHoweCRwRV7DJmfxcEo0
JlBH90O58IKyzz4GKwfCd1Qdc7MG6B6Qw27l38bGgcCYMugJGaDh0OmcMjbFhno1Y/PG1XRnblRy
lofEAp4gDmDA/02se/CY/asr97OTAxrsYFCm87HFALsJRApL4DjRS5kwi5tuk4hpbra4sJLkHo5r
iNYQqeFpidwhLINGz4MiQcm7N8CSJLhW39zAUfT1C3VH9d1NidIRsK6YkrZkgjaxGV8yczkvCwqg
AKhdly1bAz8hPz4BJ0mZSurHe/6PJMTqEn0ErDTQ5WqjTYRJaKAGSnppJ+Vs5CtfLp3ZkSSo8OnU
KrdpPElULP8k6DyA9hiE0PBrMkXZFdjh97gLIYmi7rVA6w8qlEv7j6qFFj0ZDCaxi/CYAcLDNSmd
8KkYOhZdNP2RhJ4TWo8RSdfr6h2u3EqJAvxrf7ZQ2NO+bY3X8H457AObW1LGA30wOYW+y2vftQt4
Ji0rf2aLu4dmmGhbrFA1AQT/6fgSqvYfOK6JSc03vrOjuVSFKtkQ1xG8jrHXHe+l73Y9D0S0ttgZ
JVGVi4j2Bh0vECLBe1wzI0jZbD9g9qkSEJF1DQ9W3pUR7p2Um82Q1TdkoD9wuTJJ59NL16Q9pimj
GVEu12V84FRT50x5PwOmZSx1axunzSHBwjidDjS5WhHRdQ5FQV9VNpv++mWNzTZIkxqowLbPf/h/
uyDcrmUbadDIrFQrQw9ZrrMN9ZXdT1D+aMMBbUyZ73AiiDwQZ+0W0ujFOhtMfeqcseFt22Q8y0L8
B+wbuAJI5CJPOMHhU47NGzA9LEHmh/AoP33pbFeFbD6uofB1LzDZ+9Xy8wTiGCADBFy8cH5H7qJR
/KAarZcBMhOnZ9y5ShY7wjz7mM/+jc+ctAT/S+ZAEcd6ZU3KtEOyKpu89rFd/QadS0mJjR4zfdZj
tBL236/HJ0B4m65WPaq7F5q0FW+eraupKD8B5oJLMCjp3632GLjYoAKJqdPW8iN9g1C1fg1zE/R7
sapopc6er9aZJh4mMjKmuTTXlUXGgjc25A1TdgYCJf155YiU+fwoVTJwtZxOxh5Btnjrw5ZBuqF0
RadziYw3zpmnJywVS5EgOEzfEmKQ9WTtrn+GzcqHquIQ7ppiUU+Xeuhr5sWyW8n7HtGHdVDOrITL
DPMt1xJcilCGmDaHEvTmQLMZhTZtOBmxIGERQWtGjoYXm2F1HYlmLqne6MeX/R5fgGIUuYC4vZQg
nbjduwgKSZ6WENgDOmZQM1ZkRju5dmH4ObJPD2EgGglsHuS8IH0voK1wLm0xIOYwc6FyoMaO7ViR
GFsg2mejXWydgDQZagEv3uzZxCQ94ajT7SAPt4flzqZSnnhCTshwvEqnD2WdETcGpqh4miHPYrGc
PgYrNMQrZxFq3R9c1OrxjHlFUy0ZjJdCC9VIQAVg+4Rg+GojhBU2keOrh21GqvSxQAs3Gt7kJPi7
a4qwN3nPn3T9TuwtXdkAXqUh27Y4VSL0dUytw86ObTNoLFXOl3Mo9Td3nL7U0wcefsX69k3ewkp+
OA8+YHkTV36EeVmdYc/AqeQS7M5UmyVSQcoO0ch7rEMuWZHUdE+66lkoc85hLIvnQ/JjJ4KIl/74
mdexV6V3JQ+7CDAt6QxSf8fMGMbQ072fkOt/fma1PBwpU+L9Q2MfWBxO7E5iUl1HaZxYsnhIdu03
/upaJf6CuIx1Bbj5qdS/BbYKJQhPrSvui9do+Fvi4KsTiVYv/qnxR6U8ogtx3KR7ivDkTKsdtPqr
SOYD39dyYaovyVVrES96tN9w+BstHIWBUDv9kwxQZt1IqX0BB7iCowZga8REQ+Y+3pN9KgNZVw1S
9gyGsBgzCmEbfHfGj8sdDrgv1HUW1qN29DExTgfKJQ6v/4M0FZYfoo8/MnM7R5zQOSkWNnkdoZ2G
U01hPrTo7rHqbEJUjkUdNZADX0ffCP75u6P4ZoN7dCXgaVXJfqx87WxAgXKf9RZBwPbOOp7XsDU2
t85osf3jUmNjk+hu6xEgmbZd3MOpt4KiaWtHcfoyFSIF/dh9kjH7rwehFqhS5Cqe9+6PXvQ7+QSU
WpoPpKQy9H+S+lNQSIatf+pKKjro8hRzaV9pB5NE0n+1nNiN1NKM3B6n7HJsF0yyIxJQ15bCEesV
iakrqx8vQD8HfJtXqO7ovZ0QMaR+gai18rMwbzQJsidLBUsDA5Jhn1pw3ZG2fjyGpvZdtR0tK4gH
jVjtG/16+xLDENm7jLracGdKixuPCk8QzopWs7wFdhmWPuApRuI7ng9vONoGVPHKuyyIKE65rw4p
zKS7M/L1xU7TpBp0JTjdwTOLP+PkQpeMML/K3BsV5BdafjccpJXymszclY2HwhUgWG1qZ2k2kRuZ
bHL9pT6QAt937TjWOCMcCVASh7FeukBYtKLR1SQr7S70bV4X2Z3BQ9uRpwdD0IZzgX2hyH7QvpPl
I8xwM+6+Bp+v+KIFt+WDoRaR5jts/IzCLoGgLKRBrC6CtQsC1ihyu2gg2z30VhASHVhFAwhO+kGq
qVDuB9IpKDzjuZIsb0kvtKqEP7c7puC5ImrCKgIln16dIjyGAiAW+UU0o8SEXcXGVnpSA8O1BojW
osMpQEMxWtxOqpNevxhVm89mVsOWk1QigdRDZWn67O8PoE8Ox6crYlv/Zd8XJWpK1SucVzY1s/bo
JrTdeIyKHoF+zVvsmjpuGYvjjkWoHTi7PxZf8MGgD775QsWvEzkswbDtVF7Gh9TtZ2Bs+gD1W74Q
C06xhDTTA3nTQde0WXqvslXjjZEnLr0jyqiv/SwKsRlD2/9IW5HXAK+ej33FOPnNuuwkIHxRf2z5
8fFIo0BYttp4h6ThXm44qa6pZyzPJGpRm8/fLAEEI6gT2yUbHzKyxXsIauSmTdswYLy800029eaB
GgYDQy5+rd+c0c4jGPqBXMeR1SdUE7OIxdC8w2kgJInahLkHsWnPsg9OArXydU6sNJbIa6j2hZat
e3u9b9c1dGNh03Ujndzpvi86lCXiF7xkiRsPuXcWtMfIPTv1KcxdUpWDa42OsBc8p9eY5vDabaqm
65gAq7CCY6HX2OIsZy9ZEPD8/lCEKozKAiapIlWP5oDib7aAjwgR6ZySp50+0M3Fc2LVyIttefjG
0EgAfHSLo8a81euAnL4c5Kjvkya4/0bgkmmR/j6itWZEV07DQZNTYWWMST1cGFP79qs8MZiH5FeL
/Ls2ESE0ZPCORsB6mYHFz0eUAz1K1MgWHScrVEy/eoUh7PGQfgdrcgIsX1hlw2YfCLcb1wp4bIWz
CMRBYQkPc+1QeYVd1cxgWot+Frxpd9/JabJll+U3+vg97bHgLldScF/XRFz6KH884AT5ZT9H0c+b
t2w1RyPWroUblKUXJVdbivl6Qk/XvkwPiz6mPHKyLuCcNGY7Ez4n7JKilzbCtND1V/yHRmYZlOQu
nX+BGJW0f9B+CP8zFg+sIpxTRYZ9wI8BOJKBiDjnwfaXFGuK5vp7EFJi9mSG01WKtMggLWWFiz1N
729l208jXaVotThqQPRrccf5iiTWrjjadRa2ytdiUKXQp0/b13cbblPPheDQapaZfM3X5hkLOYQv
Gm5jiQ4keE5TPoMaZLqCZh6VyuNFvFtNtvcueYp3BrC04fWeM2Ffcx7MdytCttzjThfs0FcXjvKh
gLoVTUZmfMUza3KP9bjn1q3cG8KbcpAwTyKpOTh2injOSGz0DC+O3cXU6VQcoCnlOLufrM+TCkbf
Urly9qkMHXQf2ChAh7bGh07EgEh8jUihg3w2U0I0jc7EX+cl/7Sisbxuq9cgV/a/BqnNdYXm7z9m
0uiabadrQnX0VJH5oFSsvWvKUMKTcEnucHVojxbHkke4XM6Bz9OfcBObOG89ow8ur0vUHpciRf/S
vZvngkgnQK7WHWRTrQfwPeT0IKT06dsH3U7R9XmKPY/QZFNYm74tClBu0EsfAD1P7xzM3EQgIr3H
7NWosE/aQga+CmMoacK/3ngL9eT8oN1aRR1AD+rXbC3r1vdU5PBWmfPgSV1niU06qed26QClgJE0
h6RufPsrWB+3tPxeZmwgZ98hYQF/yFcGhtQqV01QbyMJ/k73BJdg425yMdDjsBF7i4lJeeWmd6KJ
dUf6x9Cf1+P3IFCorOJTuIy3d2LNuYo/4T2QwlWS5EB6xjZwae7A1EBHBJ+kJhA39BHzzz4XUzhd
vN6+tSRlBYPI2U4ueD6BhLtsNAdunXTBEPuUIrNZh5omVWRDOoOtz02ZHoQOZMTEi2UN95cqWwU4
slCOpvzX3I70ZqilvAkfXcCUiebmZk55wZs10SDOYma/fgEnXD33ZHUvluhQoyhDH48UGrRYFrpD
eF2/mWmJ5nnT77ybqa7GI3HAxMnauG5nZvtCUld75YxOw3xXabIf6e4TgRsAhr2dXD2nI9oySUi9
OG5yHS9xInjRudsvcHYVgeRv88fchoS49/CEndF0krl6udOEY7f22MZUgnG7BONhPHWLcquUoX3B
BP6ybEGZlEikxMncEJ8u2WDhuAxl20Tz8pCFBiEftY4vS7blM9YeIdXzotG2/v9q0cRvYUz5JUl8
Nj8nbv6gJfaGvieGWF3JRwNm55PBhJ0VBVcxDCwro36gpctVOVPW1OASVU04LxRweO+srerxnpFm
MhPx/jwpq9O0EY3JMuxvFBA8uvZ/UDbP3RvXsDjiaRj0Hmbsa943yG2zj2LNi4GAukEGntnHyy6o
FeFhRWgI9tjPb3yIFeMC7uI1udjnXmKQpJDDcLvqSxVnRPdf+IhiNXnogdYijc+EOxJaRTCJ+3OO
27OpkKHluMFAsVV+8r36mDYSkNYLNQY/ks5GcqgERTN09gWGhP1Kq3yevgiU/iiOCGo+ZAkENJX9
VSXaRy+SGcgHpWNWMVhGO9hMA3CKifzMpoDf0jN+6c/3sBGFRg9SuoGb+hLuoEM320tNbgaKdDAX
4aQktliIii1Ra1A6/cHhlF16uexyYkqthH6VA4XLMoqo02WbwZTV8UtCyZCtAWVSIeJj3KHSnlKs
RHW7iQb9kDNb/CxundetKV5wiQ0yYz3cimcB9nsA+y18WnRbcRYvY8ArjIgaSNWCJlgub03ITVnZ
yRduXEdxrMvFvvl+KpNz1RvV0eGveDKyMYHQuxnv3XJnu6KnWeIC9ksrdaspnqakqg9AhUvFz7li
oD8DpgA2Tbav6q6ZHqyMdZtfhaTt1CCstM5txiIOQdUUdiLrLOcVopbSywOQhgwSZxeKrJB349sy
g0J7I8reGeJnsuJSe7qy0UsaQogqlSAdmzAWxh+b1mmJji15CJIkpD5TGd1P6D0KBqdJZZuMyx7q
hJlxsWMYVnUudt6FzX0isioFBYRnu5zrOkFmDQI0GfswIfE+FfwpE9SpAESEpJoVKOpIKvFLXOak
aecjnUR4y0r1z3hXps2Awe6pRTybE5f+cOqwWkCxdCWjXKQJJcyKTgU5EFLIT4CqiWuMinHvQdjG
AcZqMGeVb6tR+gM5kv7fMNFVYwaSmHNwtOmmdbu54Fd4louQ8UWk3spzO25hnX0GbUrCMTPuPmnz
bNg6t+HpS0Iq+5kvVtIqJtUtO6s7HDsq3EUVfMZTudxZR1sKpiVBjZW6WDYsZEhkmJ0ztnFgKotm
ttMyqeqaHH+NzLusXEryd/RgjHzGiGPZVUkUB1m7PIDIIyQnWTFSHoXS0XY7iA1AfBz3QmarozlV
RctOZxYgmI2hKwTjCVM1kjr2rV1jFfcy+MYPMW/W3M1BcV2PEz2fjQVOztqDjdCc8N58FEGraxfT
Ngqs33KrY8/p7WoOEwQsTNhnw9XroYG6rjfDXKgkPBKr+h8ygUPXVamYvaSJ/czogWf9ytPx57gI
64IjQulprjnbzdI88DH3uSoJ5KBngdCDgit77L4UG0f8pZKXT2eNBibqrPrakqEscfXmYiHEZ7yf
T12pwkEPeXtrYyKPljKjXFRu3V7isVM3DaA5D99b2vV9KM5g8pM69l8nzE0HFHfwZ5qG8WbyQ7zP
S+fiV0KriV8YHEcqcgBhHbj0Q5hDI+AboWrQxNe3bpyGGPfPme+CQ3Odbh0ChnbdU6E0Ef+whGFJ
ijhwjSR7SPWsoGkpG4ciSlHWSz3cT0ANDGJIn95o8sithMo1apHvCRtt0N8d7IcuHQJgHuPCVXWQ
JngPa4KXwILN1MhHxeBq9EokFp5ZsBkvGdPUJ+5+vKbqvQkdhxNaNEmaegtdmb922xXgwqbyRr95
rzwbv6/oMLjGFG/nY3tExriPodfXj+Zx38xsPZCchdpob2eLpZNfUA2P6gFNeXihjI2W0i/5yLwp
sIsNKj/lkN9fzgYnnLUMh9wO2Q3dJFMZOl5qB18MSVL1txTcYOaJzwcv7Bq7pvNnIpGQ2B0ivPMN
LyLCZdLX6OrzyjMjry64MEQq2U2GBtnZKWNFAmIGxuf/ZdT5CGsR34kuycLImLWzr4x18PylJJmV
b0mYZykNv5oprB+jgemppWd2fK7TBko/pDr5XAVXKk2z10TI+wu3i/La1A+YDSuyFpheNUBdM9eh
EiWq2Cida7d9I0+YzGJgIZufK0Xwiq6WVXhNMLrYq6JpP4fbL7my2zFFGCFLWtySIrA+DFa8o35r
O5IyaSzjRmCnwTnAP7ucZXZQj1DxacVDBE0t2sjifHO5ggRqmCO2CettWB4MuhMidXlPM7eoZOCR
y0lZf9gdLok4k5OLURTD+AIGQLw1S6wSjHJOcIr42nrERtdqD1zpNMGLpJQ3bC5WiomspeCrb7CL
1Ei2yUzijvPzgzY1c6eC9oLnzqHkPJ46TeBWTJVr0L1gr5MxB9wy72LSFYofgixKhywYJ7+Ea5KB
EfMJSsMHxP9qyPCEYhe/7wUGhZuBi1ewPf0O2ANzdK0xwhjlRVVF9kymRYwFay1kuOI/GDk5CXfR
BTS59yjA5teoWmBq2u7owMhjsmu6cO93Cyz8t1HAcIMcMzfVL3JyZMQb/i09hdX5wSls7R1dEyKQ
x/VUj8LgD8D3nhn2ItbxAOWKsEHwQ6skhyIq9uZhkwDLqKksyYCF8klRRJqszNCYVMXglhw953UJ
FhaMF29jweAZ/JntAkC2Vuq5r0a2y1HHKjdEhThLdwF1ojdgS4Laq7RUEmgap1AISzgakoLXHcXb
BCULxw2z8PoWQqCsq3nO/hffveLDWqeLF5T7QICmERzWN99CSOwOcAHmW6mM0XLnEa874iNikbRF
KnKGfigEZzP4Re3yYGXwUGkJMBCNenfNfGH3TUsKJs7Bzm++7e5eGtHL2g/ZJOVVrAKlopSmVS0n
smikTNTvEMVTbZcSKy3B0Twg7Ekw9fIpwIB1MWkOv0K6MfLc4L9zg0AkJLXcKBZCh1c2Jf6IpHIz
r/xTatX4vTcqgIT51OpimF2drDS+XBL24rUaOJkIBPaK9ueDrdcIt7NcChjjuw2G11Nqrqs+dhQL
q6LccClL9kytoatTgXfgAfrOgkqwc+ulZXrB0hOpJn8Ow4DWsfb6r/XJvU0I6NG82jlhkux9fkUz
KqOV5ziJvIyKgCrTphLKadrsEIrKt2UULPryOezhSqxfl6VcWRVyaKByuoDsGSjddDIYYwenayQJ
TBn9kw3b/Lp69GOYj0QgCjJP2cftBcBTuKEzW6Mo+oAo3FiZA80I6IoHUA3vAbsGZiAfvRbS4lGo
0ogkUn9FmOqGYT35bDkmM+7i/Nmb/A7YTLxlKw2tSM/QKIRdzEB/rfT5w42Oj0eky4LubyLU8ifg
59KEHLuhaO/MaXGi/NH1xU8VvUIvbd4MwQVmAmQm56Mk32rtoWH2gjYpXOAU+TjSGrG+iHEJyooy
hKzt9O3U23o4Ii7baV4MA098OpVTACZ9P3q3Vsd13NPCbTU4cpr9lADu9moxgXVcsQ1WIOKhHG1E
rEZQy6SMPTiud0RlwRewE7W1cwl4E+vvvlxU947SOmEpx21Zm4Pj2ZSQuwdNUnUs8km7s5WfQuhN
VXIzpCPJS9qTJiAqKIeZ5bwx75yVADMHobJa93yO5qzbxL7nC9k/FbHBWgsUIXvfUWAYJs/UEFmd
1VERsZqTzjd7XEvSZedE/fZDApfDXdKW2nEqfU4yfJs+WC3IjnhBUdwzaz6uXPFyUgn0nHci6Vhc
mllbpDxpJT1hAZqrqgjMPWJuJ1cCDEgshCPXtaajVxaEiEzJ+3ietRCzaxqWrUix4OV33uW0Ke6x
aN/hYpeEf8r8I8/8qbL58V3DxLQ2AyXzAtwfsGuAcgpdUWc7/UNVb3rW0K6bUeLJvi/6WL5IMlzM
gm8B9n9GJ1pSn9GZLIu3THAhrxC88c1AE6jmwvtkRZtY98DR6EBqqiLYo8zxs580A2mZ+ww73tPz
0XdsJy72IwzAv91XO9f+lRlT4PODCyjOGaqtlvbFpgyPMqrafxy9VD5TZCHMC62T7xHpXz1WW3Ce
m5dl5g6e7XAn+7/ZFuauYsbhcm1nPVDG2HhSWC2fr+HHtdbAbvgr3HqW/mgEGVzvQmPytJSAVfOD
f7KCHn9wycDN00LAvwrsl+zTxK3GybCn7ZaLfvK87SOShTEUrlgz75u0cA5mI8B1NGDlx5vMqDUk
UL+OnlCREF8mGVb32SRZWalv89CtOKGOZHjlNOMsdUVo4d115tpe2uzbtHN4kRJpqAlrKWaAfPjz
rzuGfPp5nBAsVz2ZcP6M0ohgsUZGavTzzdPG2ZHnKhgth+9u3dILHxCnEHVijyu6jcA2I5G2LMYl
VpuhCpwx4deMDCPsgSB1UkNB/Va2CtR4WjX4Y4Fo5hPV3O2fa2xNaIC8ZCySiXM63xH5pJSxOHfD
gayN/9JDSwkbyeuUO4MgNToQqDEx3hMVAPLLRxRs3XPc2ClJRHgz/7LYlIBqNViMDqyTRiwFviaZ
emgU23e/ehDoKu0/6KSGoT4tjhRRWIdxwQ9KBc3TQ3kmjJpXTcPoj8UAdWN3L+mR6DuzdlkVnpwP
k7mMk9yh7aVI8ZTBS6uSYvLK85NcZvDFnjk21qPapWbnWKFUEG5wx7FLny/aSsBdGZUnIpSUHF+X
+D3kkvq9h7AEbeLMKp4n5NfXLMmfjgh6nyhFmjY45RN68zHaxvVtuTl74mQvNFI3bebax5qF00z7
ULDU+MMs7EWS6HZnv+jsG6k77fD/XWyzZUEoWUN3ZrN6E0zLGZGv0qRYheIbHY+4hJRHgBYauyAk
/7Z/7srbDXcSX5HVVYtVAEBPdyDKyplDqRKAiEN2wUsHI8HXc8TaATrjEPIB2YOcmBNhL6DvX00v
O3jBlMUsEFHyIjlQSg0v9GMAiALETOcKsYwuwbLO7tnWa8Feo02VGfHMcoBmAJX2Sxput9T/6zDS
JPSW5nHRX8GlE/VfsaB/XXhXuXLgRPIxAlI4Ram/joqJtapqMS/jy9Xsj+n6QyI1ZzYMzSr9Sq0f
aHUmZWHGK7nTi7rJk/p/vPCpgqOr+1g3BMAAgamfd2pv180Tzm2Xwz8tK60Qog46B7X533+kaKz0
xNao5wX4aJMF4/qo/GfVICj7fzpJN6+d+YmT407v4Aa7tzluhvzNLzifYpZkfQfK9HDfGnEh3AV1
5332Z06q8Pp/X9PHqUvlk1H3yWQWNHPmTGSvW3aA/zrti/0k1/m5tyDjuLaazjM/DVJG6T+sjkmg
496w47RHP7spmJBeFnkRVR+WI1pVfgLlG1mHgQLKoqF+wWIl7Y2/YUyYunXocpNe9q8D3rQI0GlA
Y8MfT+3Oyn2I+lVQjDWeWGDxOcluCx4CErVzttNm22ZqneXw8+S7kQJP0T/3eb1mowamU72u0osj
cp2ocCBMij8aZXwt9oKjW898v84NdAGjbAU9PQHFBKoj774qySSIwtEA14aC9fkepV7uL0gcFtG9
4KO3SLa0zMxmdNFy5EPXGsikE40a5olrf9bgb2iLt0A8T97It65lXeW57jLE6L7BLOGmi4dOya6I
k5HODmdFZ1EY4fvDckIL7nPbrCAFcFM8XbT/NSh3QLIfcCuV+1ERmajJJgvJQRGDAU4uiY5upN5B
z3Uy5T12r219E9SyqCvpoFq8eiwrKpZKLT73j3s/nXiSL8W+ZTbD2dPC2hEoWICFDsTYIvT1D/qf
hEttAcbGUY4Jv0gZ9AII6IgI+qcUsyxnF7tutBfrFte/YONYgwvrvA0LqLZeLRVKXuu6ihkk+8WR
vWkt745ALda7Wc/DWIomn3B/C0+JScITiCJ7mEiziTljmpgeVNJO3DVDiskNuu6qEToo94bGG+5Y
Ezk2YrDvl0mjwE+fCWGDc96RT93i8CFMRPAjBh/GDvi21FFt/irPv1AqgQ9qAA5VVsNAnDabyY3l
ed43LGmu5IfPHnErPfdAcpIMCL+ll1Mw1NjtfL/B/JGYV7U5OVG5E82lqS7tjh6c4rf1Jr5/h9WP
2hAGONM1op4xsmZ2v09bn918fhw2qkjCg/8PNbUB117i+CHMI4xq9KXKrmsVMenJKDUvWsm6Q9Tm
58AzVmNkd0Od7N/y5cSXyWCQhv1At0z+vTg7L2SztAhMWobGR9U7ZZMAboxW0uEnFWCSJ55LFgXL
5rnrJgIXndIw0Jt/uFiFKE3QD0O+yBzxc2gHHcH/ppcOs+Lk+Wn2lBUHwDGx/yTHgIzVtSSnufuW
WMSdZirtrwAlVVjcKgH/nx5lZvC6FzPxTAuYh1WCsyWWaKru2FxhiDY/ixa++Wxr+3I4JCGbY8tr
ZrxK4t+IWUI11kRU95H0Fggyi/v/0r8G4G1xJ5HLTcWwVeqiaPhicXujW8XEUOuaEIGGGcfF/R3v
i/2Csjr7c1uyreQWcobRd678V3OB4sYjHjhXrunCoSZL9RSwWY6CYYp5oTXzKR+Tmp8h+8/F43OW
rbNfhGi1aIv2vsfCcrltaexaFak/mZkdOWI37Mu/VLNOrMWwk4AFXMsS+tTv6tDweonheaP1R0vo
Gtf22ONBJrHTKBM3Ch5txL1R9rZdzD0C77impFpfA2btfd9c9HS9XU4mNwZPEdp3eulqcBQ26aqD
4L1Vm4NqNAcMcciOluz8vMtQwTixqcT8CLKXVTwfYDsh0HYpWgw53R8sYwKVNXc4sWkTW5YM9cov
8e1eycabidk+jMzVxPibSliTD+4tZkPIM6jZlSsr8smV9nVgA8hTEFxpRTOLE8IitTb/HRM1Kl/L
v2ZmuGtJ1yo/pYiUUN2ymwSRGLlcXpCaKXXgBE8520LtUqOvrwdvowqF+cW5jqACggZO5dTkMbLs
GHAb+V0A5IU0fmZAzkLo0eVhElXkB4uQQ4LgkbVNqClwOUHqXKQUQm+JyXa8717EXLmZhPKSP8GK
4o84CzxgkAA6e9pa9e5hiFhoswlf5yxVRNk4Z1QG5+iRP3XzyHAJ49AVPz7BZkmoQWuDwCblsCBc
eJRtlUdUxMn2c0q4WI60oh5HeADrSRM6yR98geV7Ho9a3S8SUHvbXbQuB7Ma1ZFX4S5rQkz/xElv
0vmgtSMSjZXOEVXjtkiVC5k5C1yQEfXQg9g/Eces8pVLLT4ugnia2q0wLL8U+HclFDU6qU6i6TBg
znFSnRe7HbkDqxnEqlyVirnIFAvBI6hSFJbhVssE8GwPSyIWhnnuHjWH4srpUnZW3H89eD0RoeIR
oKzt9T4UfopSPjuUJs60edfV/DqFAKLIBpvi64quEcXr5sJX6RwRavvgsEfPGmZRbFDabzUXbhDA
2x55nygoy9Y+9qBBC3mxgZGl5odQzEMRs22lbK69YXpt8DNJCTklMGOdygKJ89+ptNRiFCpJYYFu
YqmjaVtrz62DvboiZlEtAq0mz4vzwg3lNxwnGLxTOHryjgY+AbpelVFOgf8s2KzWKqLG1W21JZy8
u06cUiBb4TuYHN6/Ojgqof9oJcQRMuGdI5Fpcim9Yd1zIU6TxNkC0/Z6Qg4ngQarb2HFtDFOU3qs
lDmP+7K7qoe6UxtbxrArIV6AWsqSfNcfTsTCXewOBUBakfKmk9kW+Nf1nvMoNWYl0gQt2kP0rGBQ
m6HBNGyvNN+J9H8PhaB747EPqGuWI7KNaS7+dWUjIIVVHMYVaQQoNvetd8c2SQhHCSbjVIzmTml4
taYPv1f3kvhjeAg58PYg4Hhc3P4lrDihY9CwxFXmhZKITOvww2ZTA2UX6fRv3YTSVXS4fNMO3/Zg
zKloQswaXTjQzRDE7lc79qet3BpVTRYe0qpBYrgVNjSpl4UsK6EyOLsjPZqoQUhEW+RiTBdCew7T
kM2Ub5q5rm8WJoxcss9om58faJE33zzDJlbFymgVuJZEC7xtc5Do9fIB6Po47elojxgGOSXwxTpo
esouvgaIPAKQTPFs4gecLWHPOEWwg/qb/E9jju/bw+odjWOY5WCJ0D/SVI2p+rWWIJcmM5pVUoDU
8uN7jegOFey2i8fsLfGzN3m8xNZNrKRmcqKqXSm0MHXgc5cvv4KGCxgD5N3LsPLiDLDPMcNtSDzm
4kHQBKJc6m8rnTJeJaXv9QLLJdeGWyLmWWuy9veNt5h02ZLEDQlE4JeZ0CY6FVouGqlzd8tqT05u
PbhCvodFwD2oGMCIKIuAQWffDkRmziD1ajJKj7ujbsxnHy8No1XKuyykT/YCP34lQ3o2/ZQln0X1
RY0NJq2Ex7AHHOrmNd/thOHyIOPPAzKhfTd5nve57vY7E3Xfz14PAafC92A8lsYJma3Zy0rYvWY3
pvzFNVwHVzs79+FbfKNpwRvkVwpl46HpxoeBd4nNLpdZLQudhAXK9vGiFRMHahYlk95y66Xwf442
+oJI9JCz0C/X8nkBZitv1Z9+i6kKXaCar9umBgpFxsIEKe2gx4Y1wZlWYQSN87k7d3IPGwxrOAzl
9D2jDOriH8jYYfMrUbgJgHmzXtfbsbjiNibgKiOOf4IoYVWyDE5aEHLPjMJ6hAXmdiohYPc0Qbdc
S8ouEO5s3xj6By2o+IWXHXOmFh+emWBhX0G4OeFCDDzQ48pJV/YY6cQLVLvBRe3OfkArQU+7qZTI
HZ/JswY/iUSzcKp2kNqbpqRRED4MiT/P08ztADuTiH8Lc1C1ZsA1ZTUKMBgcIMv6fyStqoOi4cW5
S3TKr4Mt0V3GXilmSAtAne1wWuW/ciEzWb7+gsWtHMPZV5inOWJyg9H/deOiJlJaUHLhZXsHZPx4
zOeAmdHnFrVm6gJiVbs7PgjPuDGvHUZtDQidtSoKK/IGBXYX3u9Lk4wdx2OI0Xb8Tc1OPN45NVgX
767A7B4MrNEJi+u/BOjuTBoNExwTrwu1DYwQQiZkV8WMiONXrW1C1ZedX8T2poiyGbL4zbaiu3Js
td36G2Jzx3D5SMG9N6HLxWAohEjBPT2//eM1xto4+41HI3DNup7tl9nMT2uNcfCmg6d6Vv5d65sY
lHxzm521VJUwRc9cVe3gceA78LwaSnNlZpBLCyO+Rss/nJdRPcvotbDir04aZweUmJS3VcWAol6L
EXeQAP0rq12zYWpPyyFudenUNbhJHqgf47vciIruuxN/fhyypXWeUzpjjY/urfpjhFfttlIZcCzT
vr/m/U6pA17EJcWchPFmL0UJ31VL7vZGlZf/liLhTeNMEwPDg7fAKVKqit8XovToCTezYAYaRn+O
2F7RgufXXASz8eEwonrrFXjeLBJH7bYgceUV/2Zu9wYRZp3NXj1xxCgFU9C0qWbG03g6l0IjMsP3
o6h6MPLns6ShSogHZ8J8+8iszpWEFDBWi7PL1LMD4seGPzgKPxGTbriC7yXqOQSsUgXhvaSF6Pts
fpEH+rQXR+Z2C2LPLyQtcwBOxLCpkpEYnncv+OtokM0+ERvvc9oJJBfj/qLopXr4WjA3AzzFlUwY
h2FN8ZA/keSaReSUiNrLxTzDcUOSOlbVHjxWjdBsNxhAA0VAxboGa6RN2VgfV5AyZTb8txXHtQA1
CUk3Q4V4rWa0tDr9FvNR5HSzFY2NCk9f0yLmyj2KCynkSwrIYJwdW3OEb6BU2dAuuBkiwrbADD1f
wd/QDK6PzqRW96wGGjtqHNlm9XIxkYqKIDpXG1nwiv69NluCZOQLgwJnfOy0VG5KDwDDKvnU9nT6
TtB/j0/NCn9sx+vZkkw5EVVQCVFjzJHcCil3dWd/GDZeNMJvpH9XFFEs2CK/qI2sLm3lmmpvhE0F
zwAhj06WPRHARlb5a1lsmOeozzahfOtf8Kw9r13HJivk+Z2Q5fpzfvDwQu73ulrHYjnktw7UZZ5E
OhiFNwkJrZVsFCi5+lGymDtxq3Pvj8WWm8GfS8LbAdPBfTqU46iYL2p02EQ4REnpoPYnl/70xPDi
8pdPUdmiUNRv1CZveNheohj5p+LLcx8GerX1tbX4A4EjmzxXFscET90lzytiyCGkBHCVw7oQnMoU
zr7TTlwr9lN3f7sWzbxb2Q5dk/4kK9trncF7Pvszn4ZJq6Ybfo71dM/v/+yCM9zRJQ8dGOt7eLYH
7dwX5WugXuSGOTFEv/8jzY/mzn+HbpZKal/rLuQ7IvtHnbTzDz5I5vJktPFo424MfecD1Qh9Gex+
hsrofoRDz3KKIuWyYmYjD2rBfV60INKUHAesBidpa0UY8Ay/EEa3k1sPshl+7KJvETeQesuOzOJ2
hbUejSF9zlW42GOyoZhDwpeKmKer320HKOpquWFOIfxIiLBVNciB9yCdRe1RoWlQtK/wPzi54LS7
mkurI8GJ5EIKjCQnsntZE5jHXipaphDx4p5+9ZRusDEBjLChr0yTafa7LsJ6URBKh1JiCjmlyF+o
Tioip5ZEl7zMNbrIvFmVcl2a+igmT7trabPVOWv2sZ7QOQw7n8eP/oFuiIcBlxTqr9jz7QJgGM45
qeDtSwdKmY4z9IcdFqfJ8My+MP/anGj5WMzt1EIEik9AnHwyI04YXOlSru1ft/9TIfXOrCGVaFMz
AqqkwAnPaupGPc7icwv0AIAnSNIxSTvJWMIjnDhUBQMPpQ5VP1b5gqhy3CydG1yWuofTLjFdrHie
brHF+Nkt91Ck3RMdQjFqomVMQh1RdT/HuKWDlCjaP7paKxlVJRdPp14PHHmd+q0DxGWBpGa5Vz8P
Huhci8+FGv/6MNsto8QTFiUmzQtONEiXIdbq8SiOh3BkzTb7mqXJqIbXwHSCrDb7LtAOxZEFji7p
bDfpFcHPGsQXTYyG5vhXXWiLOzMFGKOxgA9LTtwqR+PV/FuZetzfndDi78OwiH5YmBXFzaplWKh6
pUCHGB9lYHNgOLm6zlFTqLQZTSdoxoHQkabc44jmgCc0kPKWFbpw65x/QNpY6InpmzDCgujaBeQi
9IJXkJ31yIdvXZe6uuk807iqlXzcOtHM4lqTj5PFvbe3xPARNOIa3/D2aDtEZ52FbbVj8bARLw28
fmYWbvvvNfrIaZRi6/6O3VprFRHzo835l7x6qBW5/6NbxpTfIceiUkgjON6ln8HfGGAQZeH24Uhu
yeHif6lsb5mElG8FKCxrW9nUhVL5jwGxw4v/P0d1+WUT4UuIOS6Nx2GoTlpjJfrv5RPb71aZSj0S
X9Ms6TTzRfWqGfdTavH2zmoR2JUv3udYL8mVUDhm1NPyjOeYuVudkaiRKMXE7o4ihnyZ52tA7axq
fe4hkbo4QoJqdYZHNzV4+Ky1RrEGg1rGYEMp/G7I5APRZC8+yMJGudAjNAPC5KXL36l2rR6xZrPH
2c8KZOmp3etxyrB78tCUZawukQz48uFPr62i9DBB1bE8QLoJfhEtXLe8krNfcu9eJ1BKx3PlPHfN
KrZkdqSLpXLEFefq8I6WFayqLQL8/wEka9V8BXHJgYoCZy+2obPHVkGlYMwoU4U6eqWl8rFR+Zkk
AHRWxDfNZZTi9CZytsdYbYRO1c+GwsdnNdi4UDI3KSVE6FLiurOrdkjOG5zK8XMT/npW/vnotZkB
hSj0DDtAXYqxf6BqehNPT9jmcGOALCKS/EcanPlip6IDHt9UzTYvPzdt/3MHeQd20RaM4uvA5Bjw
GxRVL9amamIhIzgHP0lV/e/H3X+SJJpjFHiqqKXoWCs9TjNUNnzUwl7l+C6ljdUEGgCgnCo6ZTWa
VeeH+1sEnSq3mVWhf4Q5pvCbVEGvkZuNRvpIgdlO+sdBS5L4YPYOW5kRe5joPy71SKZTcgh0P/sh
VPsJ+5AuvZYLVzyML9Pp+/Rq6GE0gb2Emipj/RSlnI6Q2luYr2Ezwxf2cSZHGKXTw5VPBNRCvNsq
f6opQnUvcrseXJBtHpkALUz6RqmNK0lP/zHsWGKdHpX+QToDDFj21nZL3EUZCKGdwf72ReaDZa6Y
ByhkDrG0QsXTD5WiTqrgWrYirqTWKzu5NzReDfu55cQ/BBxE7Lsa5FM+a0B6IhEMmyL9+dYvMONQ
jC0oCdFSC47RACe/r15lMLPHJsvfOSlWz3g+zN5LjXHSKL3SvOgLx38fRGuiYEwnT5yLnGlAp55S
zZcOYNpZM1AOr1jnq/b8HTQag01GOXkXHLeDVIySo1ALCVIqhE6UYW0o2WMHyfq76zNEUexC87os
aVeP31qLC0EvybcHhWsBz/gBkdC1BwL1BLbCSsJuA8U2kQMnTFMb5zTQA7aMzbHorOPvkvTsr0ez
GPVtj7rKJAEGZV/yK8RitCEj8wowpAS2PZkQUn53obzI6FANlqqKZ5bLKODcs6KlCObs2BzY3z/L
BJ44jANGK4+/LQpaHYBBk3397QEm4VzKBfdJFD+BqNAYgAFvhK2V/fEx3QtlBcuDicZ3ZOZfpFYZ
c+oZUgZ35kNn7G6QR4adQnmtHSssoLjNlrFzgR3Pwld3Y+sCQB9LGzUJZjJwpUHqpcJDZchOw++l
qOzhp1CuMtKTmUUyIkbXYbZiR30ST7Ge9rD/WR47WGqQv4QckGurN70lux4Siwag93ZgstZXVM7w
fF4phLt5shvWBz7yyYFZVrHHFxBP6Ew1pfpuGOyJM2j7hv8XMY5BH0wT9P0lReyAA1hwbm/qLwcR
RonX/DFc9hpJySartL7AdxSPh52SvSfxNV2/yqeTUWXoANTLrIy+OKCthMjL8/JLWn+d1+wvXUcp
I3qeoTsbMPmUt1kspPf4ePD0DFsHrIWD82FBS2uoCJsp9N1xVGdCFtfkTpYPWMmDDP212nJqI0ew
CLpu7UaNMKUIviMbXe7oen61BXp8QSUji19pCgOmKfkQDEBCnlOevoA5/c3/FPEoVs234pmI6lez
2KEZbamUwUA3/oUKu4S9w1zelERLa3XQtd01I4SIw0Y48cVqF+/JLcRzwcTQ4QDUrP5J9ZzCy/+4
S0m2bLJI+wWzqWjgZA39nBvw4uskksb5QoB3kzJ5oPKW+7HjVajfBb/CUvd3PluWGUg5M/A+zqkS
Zl6thMPRbAPZBIhI6R3+AAwQQlzIc0wRwHd47IJrHpKzPdCU2ACUejGuasdO7b/+s33IB1xoinmF
hc6YM2Kj+Ft1TXPH8DqKSSEdDnRXHcyVoUOE/GuLgkB4+n2I2wKrQyH+nH3DRBTz/u5wb8qCIzVd
lWw7h7ESk7tMQ3rJGrB/HGea17LhNpTanqSS9K9FvmzV0/gWS31+KkQfAISn+wfJrlaY7pD3gp3g
kPF2sjedM/1jBLIKmh58EZLBpwvM0PCGJij0BKuX3YqfBu8qhZd8ZsIzmWWawUHJtsJbo+27eWjg
I7G/5DI6/w3sDVl1JjwVs+Ud1euYG6HH46jqcbaI/LCdXZd7M8YVPukeftIcRaRArD5yTfvLLUi2
r5AD6lqsU9pHUmXoTSsFtA7LTUv51FWgoPOJDHwl6/MrV2LDd9EkjnvHi/L9ZCFnO4jSIu6a9KU7
jByS+ELuLpyE6q6BKarsJYdds49D+LEQD1nKIfV2KYxAyMQcKb+ni1E9ivOxky2P+0FpUnhzNTvq
Z2c22mvbeQsvBMcg/XUYkc9rEYY9YzyuDZCSTXcNhsvUEVNCl7yh1nWqjWkDM0cgRSKMEscSmt5s
jy7we5V1kClGL8u7mHf5shMohoO2S5sxq+jiEs6XeeqmnESkut+Y6Kw7iMeBbYgW4YdX6R6W2v7I
hOk+mlkwqDgsbRvcgTeWzguT7/0XoWDdT9/ACE0BsmfZqe4UHCylUrv0zIhSUTKFtX8Xu6gUSBL+
WBHai48f2ekFktvBPREqI0l7g417PKe+Xf4k9e6n2Y3vX1BblWk4DMsaYjxab5lT2A9kjDds9tWw
IqUa2lLBM4BBaQm7W4/1cu8EH98U5LO2G3Xk3wGTariOBni6y+pp5gfE84EoSaGUkW7xhbG6Caov
aMgWg1WrNOslms9HpBs2y9+nYW8b9HsllnxqpeQJJ2C+Phz14Mme1DAMrtfUy794ZjX6ET99WxfN
eC00Gz3fCSy3xQ80amFtWY8emQ49VurC5d8EyJR2O8M2i3SSoa50W76EK7D1poCUnZwDJ91KHrD7
rOdgUu97DV4l/B+h42itU1MZlolx7G4W9lnn55oc/24caO5JC4LCtSGtHRyFWBO8/IEPgymmLBLF
WPEc5ZKoVqg0iTbYXgvczsZ5J6Uq1IHnfBgMbKr2qqrVTTkfX5sXkd/P0UtGe7FOZCv70UFLeQPX
9w2fSn2BlhkQMeX2rrZQshmuRE0VOOiFk0P3qeaFhkAz4Aq8/oCHvLJuPOylzIXg2f+aLFWUqM3/
UZjhopRsyOYGWi4MfAoeFarsyRRI3RUROPXmLIuDzjzoL4cSldNMpMKI+3cEay9v6XrIYkp/BsKS
IK/JuJ8UVZmktDoK0f1T36bRxAp1yXNy2qAZjxtwCH8zkqsbXDDneFYgmEgWtEbBcGEdmSNFaAr+
ndFjlxYNl63pDoeY0eH+/Jp0jJUlH7IVhau+nPEtSl6YHAGEwXEfc3wzTcd9Z/DGZn5fADQnQxoB
5Fq8BIY8lQfiZkZOcC5Do1i87+Bk5sx3KPVCB858Tkyi1Xqg3w/tDBEJiMorXlsXDv+Wtf7IBeCN
h/5gTwTzN6WNf2tPZqlVgYMv4X2Rj4XPZcUIcdUaWDTyOrkkC03Y9+6DfLJPLRxzY6PkPwvkVWSB
BWde8nf/4d4zXDITzqDtiz0vS2rngaybPS6pBGoXYNsOzZSLE81LQwcQuVGCq+bLVy9Ve7FLg/OO
jfup+BNx9FbiPKHgj8nsdXTrYughMnNHyaKeeorQe854ix/FvQWpvKoj1mEPHa9L4NrSTNn3tlRI
isHrVjrFDAqDlVh6k9GBGh2PqQXnd2U7tJhdlia3uYxnhMOSqZ9WWnjaRYI8Lj6MOPulQYXZ/AT5
Dzb63T1CrurKKvqJ/ZSXTfqDJOrelHRFfsGPE643S3cCbgugyDIheZ5BBuo4bO0n2yciWlRcrEHx
WwE6d4lVpDpf9n/bT3/svw/sdsqbKoprX+6qeV88Nsh+QPxSIabSloBwcqSkxjZtf/KRgQ2xsUoN
X9cC1epDsMHoNY3uuhGgo1iht2EUtcNMIZi4MfpPXXS080YpJzbpAKwHL7dYTGc0eOfPLtzUMhfG
SLvxR0OFUI4RK/ZUIhBRe9J/g/h3urEzCE9KYkNPmansmD/CAsVdg3g05wYjTm6wAdVyLS/L/6bg
fyHFBvEpXvPFnryrkmHWG6RQDgOOWMIgwLpBNAgmI6zjhZiDRMpQX/tT/NHaifPfNFKRQxlfNzNo
zJxygdRChiwfNk7Av+kHOWkEsia+FzcAf/w9v1XKW2VMWI+C20XwrvluaWykvMT9emVGE9SKd0Cl
yPusGKrSn0HqvODt8kiv3dGN8+R79bHArdMmsdbgL4j59oVm7lij6p8ZkFKtLr2dtFP/te775xcu
zdgMWo8P1vs7pJKZLccUyh7T+8Tya4qyhfWmEFJpLo85Ww+lpMIquRGv/qWcbQy4Cxd3KGyJ1hDQ
LxhMHCQMmxmANlcapRxgax5gwAngfiWRNtxBO1vP5jXBlZGkO82F+KNNRipKNCCci+V6eg8FY1lJ
yF2Ny8tMMA2FvkZXys6hU1hdZ6oBeGfcuHBmCOKYNhf+3PEafE66rV9ahbfqbm4WDusBAl99UI6p
TTvOKk4BYMocu5F6g1ZV7vvuql0Jf1qp7sYSc070Bn4H66EQJz6T9WXflgnfD7oRHPb/ObmlI3AI
jDGoRTZbxEibq0LBOi4IQzYRIA4potOZOTttLWql+PNf9fb36GXtmXzGQnGRxmBlDlZg987hJpBo
ctJOMmzb3+IZ+XuS8+rgnxkWwwjbnRyajBhaQ5huwoceIz/zxZ6cyJqLBw5HfFSG0ry6OB72dqcN
gYw24KpqqskxvzMw0VQJ0OGVNp3nF6htp3hFQiKUhh55vSVdEEP61eevskx3sSRh+/wcJVUCfYWg
yONI+HXr5OaUJCyLMelCGWaYCLnWUiDlOCNr4SNUV6xkbDP3F6j0qELZ5wD2GpIu1kdTExFg13mJ
0oC/tnwPbcnXQ7B7UN/l3dSQajiKM/6xfW4UwVj6hChxCVtUbgoO5aisr0MBf0U1KNw+ZZTdocwb
/7PyzbpR2YP91cja8jJ3BWPECFn4Skvx1gR0L20yj+WwI07NKJW26JArSworoJsnFQNgAB7/Xstp
8roQt01IU+MgaW27iScgl1lpVU3eqIPKCWbfolhxuGozoAzWTed4BQFo3GiQrucFp0jQV++kLV8H
lZEPky1C64L1VKEhoGZ3aylwxAqlFsJudftWURf0e93qaJMl23uOGF60j+w34jArwJDAFfimdrNY
fhW7Cy8/c0BrLS2apgjY7BQtWFpvEWw4194oxRKHteyuJvG+SlAmvaV/ns2p1BzOQpewk7JJMHiF
/McftG9ViMQ9yplM3s7EFgEXAa/ZI5i3Blqkfam+fuk/xHPDCmgl7z59qTkAi19wg7ZCa+uZhXNw
zNy/uim4VeCa+cMaNzLGyYnJoSPo58ytNEXKJzfzMMzwBpeO99E5DJsJxTSgQNxoCYY53e3buoZH
clg69g6o5Klr8+xQeha3jqtIFB6e0KqSzV5ako2rxQzS4eIb9EJAwGiAOCbydnpKPGPdcK25zNTv
9L/G7JFyt/sn5qpCGpStGQowUkhkntWWf6fEZGWZ9YgPT6J+iuU6UOXA/Q4nKjXSnsqWjncaRPIY
ZdKgFB0F9uY5FQmhp+XPkQBxzOouk38nSVnCucR7DxXfy449WBFr6EHOZnIHoxHao28tC3dCn2qR
XOBLf7GOz4NTcCME2VLn0Egze9KBhYF1e9ju7pRllwYAo8BYsh5fAjTq4iprZUP8rAbsGnULtQif
WcRkhA+rIBjfWxZAEL0qi9CyydfF5mDpuCbmOGSUdtQz/izsR3IbHGB9HWejvikK9+EqBtT9B3jl
j3F3TsPtzE9GfjBUOPyHJUSKBLV+CKCjtkiHUDPNmB4AnOZ3nxXmZjytWFjJDFsS/LYq3rMcbNAB
37DvzWCq5qY9ly21B6X2h6f6gbgv3HoWYu7a05OSEuiHHYajuhSOp98S96DZ4jWlugU9cIswXCgi
bJN/o+bZ04P0M2o/WSbUXWOKVFwRrj72SW4pAzGo3bZdP8NTZMVsNdjbDDCwV/eSJbewmOkJTRx0
jV7Y9LgfpLIxu7rYBig7ZtD/4Eqc2POkZYaQHOuYqXwrHaevK0PBOX1Q8fX/Ehts5yTmbFxfqfbl
9RwbrxM2f9EAT46RZ5ax9xMjKIjtKxjgt44a2HvDgdSKNELAbDPN3ph2pQwnmhTnCrLOfS6B8NMj
ozHVX3E+e6QQRupVtnN+4XbOlgkkGQuukIixVoAjtVn9OYFBd+Bks5KttrhGOtdcdlZcw2yXhW0N
A/LezOI2jRb0y24OLiWyL/eoArl68X751NzLiNx8wlPPcNkRPvqBOkURhN695A8myg+0JIXrdu9Y
edGojS0ZwuVYnrtjqqjtvQ3rBjrRU7nb+U29aPk1oe6B7kg3s/ltiYR2gE5TAmtl2VaR3RCcnd+c
N3fSK427/uJTzS1O/ejIpZtU9vXYxwLcQIIbOwkzLJH6L715DgSlxiYWCdFDiwqq71UMse46+ind
URYcP7y4+X9J1DiF7r9MWJroKGH7irtRmlYh+Akbn2cK7Fkh99YoUB933cUrDd/Ycq61OKLE0bq3
pJ/Lc2fGlAgeIUMWTO9r1CCpRsJl6XDyUxtoRvru9c8ndRJHCK7cHjt/YzO0fvMNcC7zolDUOu6a
TfQU66Mm58lJtsP0uvZVRRoyrHakmV69QhjPKSLmTIGQwCMTfntKq6F1jdW6Xz0jicCZPGAIEpDg
3Sx52A8AgRlt3xzsDe5XfuDQLnSramULQbncnyt9USniugKAdg2q2BdmfWDLv9z05JE8A6r+Fmsi
ouvDRYr5FmtgxVEcJDtIO7Pdi5VWZ9FshWIY+vq/j5SG/oLDDPJvnOO3ShAORY3tv2vqyz6mKQlL
+bXBKmPmxNmhi4mHVbvR/86wfJKWPc37Qlz39wXRpIDjUDP7Qzprj8VLObSgwfBiTGWO9smJ0hTG
LIb8zegcl+6DLeB526FeqYfGRQW81cCugjXfs7nloLMej8wgiPSBCMVUVeyZ0pIn4nsGzVXvX6e6
pZsldTpG2Ola6dQTXKBD/wA4ievVfYgxYt3EGXm/Qac9bk7SB6nXzNmgEGlOG3bna+R3PRLryaFc
dMt1fclPs9QaxXqOHhWzhuj50fK1k+/LUaVLnzq63S8lA+oRgMP2GQPEE0aZz9YNNIRBw2i67M8+
Vzl+MYZt4USjPEnNsjhgGHMOAXI4mGw1o0rRtDAUZFsjbs0IU3uWM0QNHvyFO9ScdRPs5JgaYbxG
zB4RlZeRhYy3DuJc+C6aIhcdm8+wLcfXkSYy6gFFlz0Oxzg+v+XLwuNxn3n38TTC7ZuH7oUkSxU+
TFU2EjwmmY+BdunLNiEEXx/n5nTr1vdkruIk+3W9kBOuZFDaMeXT3z0hBbIOtEK+5H8Tl/NKtGSr
nPkCNsGQGIp/wIrnRFKixkzGy+OKM1DIL/Bg0XArsL2ta6eFzWlAlB3L/BVI5RNrBKpIA9x8Ah/S
4Qiq4zZLVKrUPEUW1+dahLyQUGljqSsWfRs+Y5lrw00Iy/c2
`pragma protect end_protected
