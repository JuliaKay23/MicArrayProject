-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
POA2pW9wqjkZRlty0cHbfsvxbYmdqsKZafCkQIqmZ5iV3E/5geb/s7j3cnWTq8M022xE14qTp2p5
kkCtm+cwSEsU9Fa9vfQZynThcV9//5ijLq1ntiN2XCob8hQXiIPPyYTy6Xirk21g+YlULoCWe/0f
TpgDAUSWBp/q3VDJsBkT+6rTrZEpnNszvf7MHNBQysTvGAFgcO+YuBI4JEE+uogWM9g4qmH2pRPX
MlNrsYZNs7P5EVv5beiRM+L7c1l3rUVXQkza3bjBTk/Hn/p71xy8jdQXhp6Kl1wrEG/6rJAnabxd
iU9vqVkVQU1AmvG9xHbd3MkkRz0N2jOWB5gQoA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5264)
`protect data_block
wDDbOmgvtZrc4wLqGoUAjGhCA5VAxUtp5gw8YZ6SIL0td5rcMJPyKdq+/cWg5b0Gk0tFOwPD3BoC
g4HaPaRdg211HaY2cYiqWViiJ+S9iFE4wCMOD+wFobKMz3vfJ/M9b0uLhQF2Nmf80bJ8rk+qURjB
VPaWA48IkLdfaae+wXWWJ42rwmRbieTidpcR2B7z22gqJ6e9HzR2GkTcHuB1wI4RNm//S+sS61DN
132my+B1mI22xVb4b0ixcG8YuJLgvBlUVvn5TadMszRdXLK/8Lp0ffhXP+iTehjKYdeIIWp0N0bt
GJrmU8UH27UCkpErb7siOzrkHIYnCWPY5OKH/qg9dZ+4U+aa5mAZotv4omhXhZxnDxdROChr8d3r
ugUrmEhAfehtOraexD4AnM0SRW1DB5YpaQPM1CpK0TxMGAXs41MDxRBbUUmaANvELKO8cJ8JUtRc
BXQ3cVpZ8KykOTR8pwIECurdn4rgIZn0ZjGPI381ijyFvrwaOuyRx+wxZ8LUuHFrBH7maVfJVbhi
wHmRCpCKE3E+jdQDzlTIpIW7qGsE4lrysTEudYnGOw7kcMT8WhCnvA7jDvw6nxSIC8UAI0SQiBJ4
DpKV6Xpi3Pi+hS+9hvN3UuaY/3iSRn0D6OChv2zbrPHwW5c7Jztqqmw6XN6ZQmKtNEF0RJVTWteA
t5sGfLRD0cS0/hwuco97wMZVspSF5x7yXQuYoDYSu9o6q71cta6c516yg86wjixj3uuEa/ivqNA6
BLKfAB3C+4sT0dT9SZmbUnwIc1E0Uo0xWKLuypGCeqh6zrt31CxIEw+qed9iJKMTUOmRsE19wD9k
ORd51jAARIhWrx0XDq69MgYqsesd9g4IZt554aMSK/h6Jcqwra+pjuA+JaQoWslN7f8FRIPlFRwQ
6TWYLCCRx17GAipej/6Vk8ehSL53wuXYaPmYs6xzL8mRAydBmlG1WAQw6lpcwcbLiropm3pXShEo
1XVGzCvJK6PiYbMQvlpNhsiTk99SFrkT2nUWdlKj559j5VxWjUOVqnuTPCF3JmEJxmo12xEL4VmT
/tifn1CAjBbeEZIJAFHzWtlR1NLbjC14yUW+4xmTcyGWdrXeD9+PzvJln75iwblirbb2RmG1O2TW
egvoz1Ay8EeDC+My52/8k83IqqoUAWobfyoJv5HjJTp8YRlNwM16u/iEuKz8i/LMIWQ/kGBI7dYD
cPSvzEYx7INhDolC0RrVZl0o3NtIVKG5rScb8yyzSSa2eCDl0o/4RAJLzhw5h/5eJw5yUZ+JZhzf
yNufjjC1zL+oovlwvV2ioQOBm3tWXXsRp03y94nCFf/5wxTFTKtzS7VaBBw5G9r4aLvd1hRn55/B
cPg5tjXvLvpbE64qaXVJl2lnRxMBYtREUGsezWqTlzsexf09Zld5KoOyRRuOMBh/wAnjSeIAwnTX
PQnwk3A5JQb1yBCGKwUMh9sNnHT3UPVfQSGuKIvqK9JS/VTG0VeDYSgMiOHI/Vja18lHhvhX0GVo
MgzI1zPbhTGr9TkNcLU2SIP4XcpEqLF8GuziJXcu9zA4EQwiEMdrUQHWRMbWG7ikejjA0At0XZ+M
rMJbbHt17IzYZlg7W7WKEThBzzWGuv/+A+5d9nneprXBbqyJQDgbjyYvuhfqw+s6a+ayIaguwFAa
jfPkcfFxFWM/dWd/i3/2S6wvjKCNk91NEWUJLXcSQCA8uKO21X2Qaqb/yHbLaduzuEFDgJLvlyBe
uJamJT16qVj/e6q9zbIxBYm4dvp2Km8skQB9XhS34vL8xdIhxmXizlph5dSwYrF7viAtmygPpAaa
6i8E+U+Wd/jPy0n+D8ArIrsaNSZL8Rtv9OZnrh9WgeVhbIIyTHCpmo30wKPMzXC5nmcFg0yRsUsq
PEOLMb4KNrfNt4KDSMsakVnVF3cfaNS7cIldANEaShpvU6nTefltqqghHdIe6BfDyZFUgGExhimd
FkfIKmUyLgfH7kXXpMevlg84QFV/Urte9CznBc/PU5o8zz/+0trKQuinZHoLh153anH0WJShf3tl
89YbfHOCrha2Nr5rKGYeKXNK9/iMIYNYEoU26JfxjfwsQjZgdCtVsInAOMJh9NCBsoJZeLHWsGkv
egpxBf6KaqPsHja2sHcpbQ8JjQOW9afmAzeQu9v8V96yBi+efmInaStfon3hpo3SWmp2gldTLmb9
ZaRwhy68qecoa1a/10PG/txA7ILWikMv7y/yUHyyLSyp1Smk+fVoztolevDD62fHmZ2qjDU9Y/pP
3q3y14lrwu4gKsFPCTZyJNFoyfS9ysHAAFSdF08AnPqGjRBzSz/boRPdqO/Om+m7IFqpTc+35F5m
cazQ4LPkPSQVnMFqPtgLkhsASVgQVJ6HgAgjJtZr5ijad43RMcqMiMAzSkSHtj6p06szQBiTir/9
fehVxwdXAA4cnmkToohZNwp5FkvWd71shjYiVW6fmBZaICz8t/hRO0KQpkOXxAv9o3nu+ZvmDopb
1DXAUJbomy8+p6jbuVfPY4U5eiJ6rSsL/vnGmF4dhf0yiAirKqcj2IAwGZMPwz9lS6iM0SrQeCzV
oFLZakXKsEoL45OC48IJ0nW5pKBYkcCtEurUKchXl4OK8dDU4UPtLMUodawCQkGY+aYirc+xNSoE
YS/F5+30VRRQUzJVjx03kSORRlyY3sXxAVIvU6fVa5JTg2Wl2WB+UXz/uVERc6ULagSxts1BnWfB
eF3NHQSekKWcddcRD3OubsR0g9gaobOVz/sjwN49zzfnEIbAY1v+0MiyuDogzQnzep6AvayyDvA1
pe39Y6Ld/BMFU4hO/SV/+wmNzgl4KLFuTlsm6DY/Py/OXUgN5m7G3rMrYCsIXezD2lkNmARbt82X
8zegcG+xWUJoA3dRLLZGwD4T8dgG+YGjKHsX/+rZulsWDw5OHzMOcq1P4bPB12/lgVS5ZiIa2MXe
lnok8gpPm4NVzcStQEmAUlkp6jo5sGkM8+UOfUOz86IbXUdLSfFzeB2N9XrkDcXfwy+ePGF6rC9i
LRXJmuZS1ZAg+kcAkZbwaUMEJ9utx7S9ljJsmoS6HDLGczJNAGwfj5fyYWdcCR+b/nrM7xhMBbxM
xX0HGPpIJrfASt/94UqY2v0eNqPCYQiqPWN60SNKwFkeeDa3bhXmBelJ0+SgaJxdisB23spxecbI
aSIz+S1bsmSBX+T0Vv0EB+Jotgt5pGNswtjQsTVsGBeZAOn82ZXmvf9USFzVOjZR8lEWxBTa5z2y
C+amzeE9NxVramMyySZ2rLaUJYFoFU768LleD5yZT8Xp5iLByFzcro2sDzOjzEaF1/P9ofNt8ogs
ERPNWbz9CjIzglIw3o+sqx1C9DDy+yD2eFo9XO1W7AmYqEZY/9QRTq7WVq7upASl/xvE/PNDJpk+
HIes5nvVSCxgt47i6erl8IG7tTkKUK9988KU6R4mIUIjtmQAGXRhi6Sr0bIS6bidCcfnznV6AhLa
VHfuUPK69OGdxAVOGgx8Stuul4S9S4G8BErbA7p5ppi61rtxPj1kz/4izUaJp/lBFgU6IHiSHgpS
IUrUjJuvppW3f5MsuxfESz1LDdGaaqFtgZDhs7XSyK8zXJJ1ysHtj3DEzt1GpjkquzFPdZlFiRXw
TSeZLFvF/RXQAYWR8LDqDhfWxNihIzBNW2aGLkjni1yF5iAD/aG/gOHzgKrqjso/tKwIU8w05gcf
YP8EqhKEV95ZXDJuSOrtEAQ7av52F+UhtqxOmtlYradYiNb6h6oorwf8FpSGh54FRB1k5l2A6EYL
/XWnou/Ptj24Mtxs8aA8YSrrZcdT8KP6nipXdHAJYWkt8wh1sBwbrYbvA3y+7mnb1sgOJi5wMZWt
cRqOwGsaf/f9PSvviJu7BGo1FhL2akw0IN31xZlnfVVlPbGMEhWkznP3gXOujilLmBlRUWjgISEo
SVRwTfFsBTpERttyFj9NXybMagl9jKFXx207Q0SGCWZKTT+R/EAQ6qwwHknHWhxbhqkIbo6c99Ln
OpIONjNLHGyY2lYgC2jU8z4xHWVmXDg6/gWoKlQ+8ok2TrTVlgYr0VqSaUNSRmUw781voA7cgLhr
pbJhyRwZ5V1nqLjcJHKd3+01O7ahjL+7MXMwyzr0CWOvqXNDJfNvpQr8IUbZRR///m6w5vt/tFpL
V54PMypxziB1OR8gl6ajJrPkMjyQQ+2f7D1YkWKeyefHvHDykZeQLEZeT/QAo18uxsJTQOvZmusK
3cFMwf8n9A9eKJvwqCnTl+fi5Jm7l+Q7fQSqltIdN+Ft6lh1p6MqTJ2BfrmSYQFQB4p1bJ+kVDuF
FEMEzNsmGd9M0/gscia8YYHQhDaBMDUOGuG1JqhPjmG80IT973zo1X7zHH0fEd8u5zjmwpUWRGAq
cMSI3SwPnN1W2O94wXJwECWgzKSIIEYvHtT71Uoswhjr7h35VBRUjTCklFGivgXOpnBqNpCvf7PQ
1o8iG7bC8VWoHllJ3pa8Fbkj8RGRR6wOzA9zELOeSalcNhg68Wzn3qKBYjQPAmbh30MtvgKuv5PY
6mCObQesQLadTrk4zD9ubOsuNH51YXzmUZG9Y++SP5shBduCCTFgNggnQKiJLD6dFvOqbDDhmdSW
z32udvbnt1D2m/dGpNZm8tp1iGcMicjAA3sXVYW1CimkbUi8cI14NcpbXnQtLfxzWiU1RZXaWFWi
b1L8q2q8JYP1I1FXf4j+fxVcC6fvSeoRdBElqfcZvMRhu5oXdE96mMTczKb8MbDgGTb2AOyMVTBg
NUxs1Kofnl8H3u6bWJadk1fivuB3LFPkw6a9/jPscfUtKr8Sgsw/cMVmAUOiftuzY/tq9zTsMM31
+YvYiZmy3Go8jASsDZw8J5byk3JiBMQvdiC3E+ckwBqmqvkXX/O1bC4QUhdz+he6w1o1v/23APTy
hI3RFHTzuy7fUnvj9jvVGXLZS7d+qoIiolk2sdI8UTlPWtd8Z1bCYa+zzmdK9Mpt8A5GHnBcjxft
Wkimas66Ym3EGXC4G+Ptrr6ZtZQnJYm7IFt1AbA5OreCUejiTwehpGYuuDHjXY0/s8u7Qcayv/JI
gDxfh4SRTULXQQOUG0ADyVwbxUp4yUxsqHtEEEakvIomr57afBdIYKazsv6B23Jn8CtBPwXmhBQE
JvCaK9N73eN/gUMSy7PIhio0qKBxvgeI/88j40vTn+dI+gFsbx3WJDWR43pMEHypBkFTPzgE/jzm
LctucOf/zPLrqp8g5GuKzieUGVFFlaQn5iPTAi86Ply65wBgPqskWpcZFsRYD24KfT69l/8pU75M
L7KIeab7saTb74j+YhO+S24Nwg/zUTgXHKkBHWo7TiSylJa8i5Bhvu10dFgX5OCFmISa5OYAiBEJ
mw6pV4i0S5IrBHdmTt+mLt32CEOPLDucU9xbWikihzCArCGQayGNzMlF/08Uk30xGH+uXb3YYeJY
8yuxu69McebJXRNrx8ozDbg9KKk4FuXiBOsz6xIWP6is9sw4bj5wIiZTA/XVWzlHVsD2chpsYBUL
pyRpQt5wLj0DTiuvCPm0mqjZ4qob5LRnqXuf85Tgtfnc90Oti9qulg2O+mxTPpPN5vw7KP3ordRe
nsPYcNonrokIGkcLm7s9jyCcidjIpnXY2ojs5GFWhgImDChDLA21ym4qTyaMd2SoTXs4vGdAvFCk
C3yIsa+6vnmI3uANG88cqlCWqtUFG+FVhPKIpnuG+W5i9pPtyYa/zwaE6xBjhwrQ2opHMXpF6oqd
MYlnFE6lXFTPcvTPWJt0YpGhU2CwbHQrqFjVqwK6aZUXwk86oEF9Cr/9a4WtaNA2c6UcQx76skrD
31957TyEVnS4cu2vnQnqo/hiiqYpLfAolWYO20UuNVQcqIXIuapohAWhSqKKH2z34m1YTVVpF+x0
mewxV4rZuWNFqooYU8YFYc0JBR8trQ7ZxcrCR57MTdQjBFJs8EyuujmNfhLZNjFNgROKoBgwsu1B
8r6DKlDGJTD5svi2KFb1XfeTDZeetCZ8HHufxFTkQak66ZH8nR6+X9Ebtl8b+I6BCQAmucV7hRA6
MD8OAVPolQWPUKUsR12HezUV2/79Wpvya2hq6/9HPOcuS1jJL6qbmszGK3JfwUUYElDNKjKftj7P
YAM298h+FswUWFuNPQge+B8ybPdQ92L0+1TN4T8JEYhQ9GKLrysfOZjwpYm8+vH1/dvRJAf719iV
a5pTiXR/+6eTEzq6wsV/w1CVeeCS4tt4EBodKueiKcB3FaLr2SLZ5nzXN3gywAwfRBxXqoNns/xW
yFb0KreKWOi8cdNq/bWjcMR2S5W6SegkuvYXh/uDViEt7TGPELMApLO9xJgrl/ql8UcB8bSvz0No
1R6Mwvf99AgPYLXxI4x9AsrUfdEjQUX55+b6XgZuZn1NP7aNeP0VEKOrcyllHsmp6NG6oeDtX6iO
1yGIa8LSgF01moANnHYAJLFLqBnEAWaS5zsk2angHzwJuGUY97OUH8KaymaPEVEup6LSAe1l375Q
jWdihMNahBRpFZX9GTjsoSWPZQS2hcYPLLad8jy1q9R7qKYy6Cj5052TuvhHkksUJ023Uf7uVTyj
zNk2tKK0nsDkcs6GlTQpqLwFknIWjMm3qydBqRJfnzN93rDxHNMFS6jUtcjSsiCUg+es6FmN7ZTT
/WOYr+KfpCa6tc1w5JTRouflnDB8t5vsiHSIWBnov0ClbQV10GDjkRASipz54LY9Vcy3mscudZFL
/XfqeEwQoTfzkbBRogK9WuLfYoaIj1rULIJLwIZkkbGhE9Ee+lRdgLZxMUjnCKvWBNAWFWSiaTIw
81Tr6KO/laXqkjlY8ebZsmXQhaBvCQJe1wGDPSoWFYkeIPLIGKgmKg/S/CWn/bVIBMvCGMMC25p3
/1tlZJDTRaKxypKFJmM5PjiscOEmMtaMWpAhR5AqeiH8r6fmWTz1a6jyx4P2MpOKJGhcmRSMfq6Z
2Snxuq/sBvsap5Qe7QO0WE+PB9g=
`protect end_protected
