// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:15 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lKOWCHmMkdy4UcUUxfQVeKDfJ0DJmVE09RMYB/Tja0VH6PSeAamLb62GdH/YaHw8
C20DldYrA2Mb1HQV/gSdf0/vZSUTr3GbgeZu0Rqa8dbvTiLSmugkh+fvmp4UrLu1
2PMlBx3DjvyEnrK2n/PHqYxHVU1A4jiX10ZAr88FMf4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17360)
MkTvAPMuivEYZO55Q3i+eiYF55bfeVPdnPcBlppNMmOgH9dozD/MPsVsSKc+PmQX
hWcm7kzutodozodgDDwaT/i9tqXgQKzeJTxwo4yBRE0GiCtggrd4HkvttXNBM4PI
xCTpVqwz9sA4SHZ8PNNylmCW9aHLVLc0H0k+mOApVambklVlqhv4v+wGQMfxqKFg
b6ze75oVmAg1Yw8DobxCS3nRvrEhEgyajIwwUkTHknvWCfhrlg4/LvmwhESoBnx6
s1GwWAQI5fGp2LTeJqNyzTrMyBuZdg/tZ9f1uwBbiJqczvpmaOZmVbkChE/2Ae5N
JA4K3DOWKHRxBBGn/IdtXY9mufJn1/Lgwk/s7OH19BCfM7vKBMqI/vv3wrAE7I/5
/sx7dZ3r32zNXO2SxNabEpim0AGBdwDIO5njEH17+kG96gdxAqYtW8kfptySJWEq
5C6SSN9IgUVs/4MqOFsZncW/HZwLxWE20m6mcwg3TIf3RXvVdvyR/hDUmIYcoTZp
nY1Nt49HYeEtsvH3b4jchk68ipy/uvzlw91u5s7bB/FoP4ItDlJ5TE1vcPrKogPM
ccHrRb6vk55hAWwHwf/IQi/1K7GaJUIXLMbK0oEsMWMVtQD6D0VAAkWQcWpNbsnq
sLKRBVo9+PegwSq53KDM+WxSB25if2+SMByl+ZOgr8k0bwhxb+tD7SXSIWsiqDST
nXG6yb7TVGOs8JyK+QROZUWw3e4BiXs/2IbGsQZ2hQmFmKOJ76Prfw/kspY7gvkF
zCSSdry/lKF5HIUz2Xzcc5mOWbv4OZITJCQ4bKWw+KlvEAJrfC2v6LH44fse5OTq
fSucwPDOvUj6AqveefvRzVP+ljMlrifAulaQXOqbPWf8M47LQfDiapvlfPW/GHVx
XTxwaOJIEc8r+wtb+ENi5JxcCe4QXr1KRMDRwoPgj4lAIOdz0a4VO9TMjEdd/vl+
5+MdeABqREp196DHSWbEXRfEBX0uNk5HP0crqOuQvqK/W5WlxA13tHg5vpGholEP
zXjUWF4lxhkqT0Hgpson9r9m/9zpmoBWclwQfG4jhGDlwhYDASe6GlvIP21lbzYW
N+EZPPuedbfzn3zvCIvRP/hPqSkZ/1I8CBO3AAR0O0mlniDEvLfCYnGN5P7PXHsO
m1HEhCCGjIZH6WCGc7M+IG0Gw7nWeAU1XU2Tqb4+0+bah2p8tRbLd2b+1hVPS3Mc
DO3KCpQnJxaBr2TXQV0fInEbT9DBYSwFH4AOHprDPdDzeE5iFvy7TUxcYK/3gYAG
T1JkFkInWqnNeGd3rP9Thudff1P/AXmoc8461pitx+jhW76i0UdUB1Txwrc8znnN
3ABbjWutlUEBZxu/pBHCFZ/6K4KJMjaWAwTEPhnHV3XeeqAoY1JjkA09EOeTXiwE
rS8AToie9mv642Xwc5rQ42/Crv2223hotED29PiU8r1E8gzjPQA9LDVI6e7FACiR
ZEMzcLpfY94NfLX3rV8jcSsvSKiYTxKwIBLUXQ/h8UwLPCB8aIAdVQvOB2m7Q4OB
Ig9aQkq6vIaqMYzV3JdoFNDssYiqFaZwwDMVU3zq03BJ1MT9vZZqXiPMXuJtnHX8
8ewu+cviCB/pxwjzMy6sRkKOXZ6lS7xJ9bhPj2G3Paf+QN0/HE+gRz9DEZEKIFsy
jYkN5RSAhOiiVBFD4thu8T66/9bfcnXXAz/30+Axhol3yylXTK46FfHIRC/Weqmt
IWmeL+Aja+n6zxUfyAMZJTIcM0tsb3ZvpWwchjywo/0GvnqWQYcWbYe4usA41jcI
VIvhNtxdx7CrmivbF2+W2G1qgRuu984YT9dm2idYk6HOH0DuMaj362+INAob1UjS
ceoY1OGS46qYzDpFp2Hahz/KTU89gsR31ycNNfO7e7e69X8tllG2sFTd8U1HOVaB
W4AdwZNVgWwzu6/hDsg9/6lB2kfevIKcLOdqO5ef+kiMAxLljfWJ2Di/tW60g6L5
4j8CZh7flLj7C4f6kBEMNX3HCl6V9urOE6Ihk1g+DfgNpFbMf6kiujcNJHV6Fb2C
TV+133Xnv4b28zYY+bp4TF0v41fRdZr4zHgWCAWbIUUcfwgjc2OiOYbwN6vbzIMx
PBTQ2cMPdiyeMEv2X90jhN6h3dZKKB8BAkxDa0r0/PIXdIu5WEPuyJmhcTl9yct4
bx2lc9i/WI42bdFUPTbQ7TxFPjoKIQ9Yjf3kn5EaAUgi6pktvJZpKGgtVGR9SwYQ
ocKT60ulGh8VOX7ycNx/1WBm0CztSefg7jXsOi+B1F+LzOgELETYduPo8phmCXB1
cZAbk9Q+aeaQJbYF7+AI6Ch5JJNLsu/XyGUyS2B5Szp+MkQn58tPcqc1MSPmA5hP
nWC10jJigYN36remXar9zSuB7FO0RO6b8OIUcGutY5EhmNsPXmPZsB+iNnirjqbr
ZnI62PrGpo6CLYhVwsBMn4YZcynhyoInbWHW9frxhObMYB1KQ6Drxn34v3y/8qkF
grwv1JsSMhajiU1+aeThpqZwQE8hu1591X+ZJsrgNQYsucJiWyzuiZkDthfkCcyP
BnnjxxrMVyQn7egyNGjJjLvcNQNy/pWZxbiQc8543TKnSqPLFFuZjmJUDDVrVECf
OQVuImJmyMHHt4iJ5HjUCebU1MznDjOTlfOAjMTjj3zgDLP/m5JFulMTZIc7pJ2p
YbLQRqXlVC6gUG1ilhZPFZpEQJzEiOUIz8XShQUF7obyYVRa/HMoEtOJAfStEDBO
SwcoT1JIP0Z9RkyLLZo5X3n3w50rTUg71qFL9OXLTx37NhtGIqT+wEmj2XuWRmo1
EqMwWHDv7eTfKF4HC6xsPZzzAqgy8LI09sGS0K1uckfI0XCXvMEWdPt6b6gFJogh
7ikwqDqxZt8kgMiYJqbf8kfu0J2JlttIez56eA67G06mD4kzHNQpJuvwq8P9mq3F
EGQorYUlXt8VO27jemrkKasPOmD7PyZymVc9sANwI32nPhgV8AzNi9ra0TNrXF+I
WlJCeW6aZcpJpyyuWw133SxVJkwpi+99HNRoocHX8mrPJxIW37Y6KnklBdiXUeTd
JL9IF8e6XVGZXGRRU7WWq+pGNi53WRufO8wVzJkktLY0yVd4g2BKlIcxjqtqbdf4
ZwL+/8Q2NKIB/pywqtDPdqmrPrzHUgSOLufbre7ttqnh6iwrSS/YIkz6EVuAr0yj
AHZV0y0RBsDN+3eSE6PgQxjP7ftEFszd9pj+GhGclW6xdDl9h30dxOmaOQsEPrfO
wUAzw9PLVg+yiHrgiAG+4+h1YPALr7sZDWU1bPXfdy3w7Q3uhQpS3fQjWUZZMz8X
rU3SE+YQi5Zjt1SrGOlG+Oo5va2d20qz1Sc+wTPd5d/UlrsQdbUQE6/hJjr/9E+s
Q1/V/Mf1eD4PujjcC6DD3l5MkhHcDdpPe4GeUoCW8O3El7yHZuH0LM3ARSPubBMP
PkyiubB91DqfnYTEeGyUjMSfQKBK7wnnXbZuduxALfNG+OCwaVOIPL0k4WYk8aFD
8VGW6wUV+2To5/YYScqdHa9hWXXDPyCwvNSYVy1h5c+MLrUgspTeIVAKJW9sxO2E
prIz7eJP6iH2zf6qr6Tlv5JDkrTSvuzTxra0Avy/IfPOIGgFkqCegzRs0RD83sz2
AtMd2HcbFwqtGIO42QMNlFiHnGZ0ccM6KYbEAnsroPtOWQ/xMyBPJ6zw/sbVssez
cD8vdvknLTKI2dxVMteHAjcSBo2aWUoHic3NimUdtOfppV3Oh5wOoCMysAHb6ZZy
8HT3AJ/p8y2TMHremdYD/r1Q47aNDN2JHskSuQwspa5RbXjHch1T7lWaFHUvekzi
8aT1jmK2igN30awNQ2mSLO+12T3bGmrXWGydnzdY1W4CT2S6/rcRmtkoqLZky9Zw
GuuDpD+Csz9dvg0At/Q7Jk8CECoKeleGZTFK9XRc1h7bO7CLRC001HTXR8iHrTgp
PNTQU7GoR3hL6S6Q7wgrQYWQXKFrxGWqHNTQ6znXIF2dDIYqNCkN+oGv4rhQgbMH
2r3KXbcsD3TBRGGz+0shCrkXOzp1wAOPIr8IL1QeY37mM5OI8G7GQ0TTea0RXPiB
hAC5HDDcxuoOL0ayAVVKlghUStkZj8ErApn+cMSEbKcokkfWozDhqUJI/1Kjp8fK
2puue2Ooo/qsx3bbzqpKwV5yPkd+etmhroiAMQcaQ1X1gIOzdHH489Mc8E81fggN
3E0u/JbR8eZWwkaJW/7AcfXQVD7KUuCrYI6YA5myaa2F3CzNZu7r9e9Q8JD5FgrM
otqjzJN6JxR1RGkpfnT3bllXj8qcuX5nFuZdvfFWEwP+YDHScFQSYX9MYPkGSYEv
CdMhMqX5wE5AMyHAvxOu5MWIK3rQgZi6fxdmMqBQFuWdncfw8AznJFUI1tanfvrd
/UfIxPMHzDCwoX7l9fdHLNNuEDRITyxFvsJ7K81i7AogtsYz2fu6fCsNUuCJE7TF
LrXEx/N8DLGSrv8wRR36esYdq04aWruuXfXv0OGg6qpDzIu8DDEhrWSU7R3QJEA1
8ooZq7UpU6NMrx9I1Mn54k58UJNN5jG8zkIHPnqhE/FqnrzSmOF6fOM6vx8Mvntw
nvsrhjI5A0p9m1HnAU/Fbvt19qy3+QNh/R3DRgTY/6lbcdGqnkOURzYvK7t7gN5f
PWR+C5cFOPk5t3PEQmi4wFLkSz39NXvnYUoo5F196NehKttAtz7DvDC6ItlwH8R1
XW0R+qqHoyFOi4pQEw6ds0vO0zNrIeDHYjeAo6QmMo/hc24Ioe6kg9J6Vvx+vij4
pFCYOHtNIN7CcGPhGhBV2kpt9umuNcjFE7KAtHuV94x9xvEpLu2fq3f8jJ3Dz+f3
zeSVt9FXsbWk9au67m+RZw6vhyD6IF5KqGnff51jU2sZVXlkbWHs1MI9G7EV+plK
NV2LocaqeaekQgQ/pE0d1ClbnrwJGBh4JIfcPCsG8d/DnSL5/zQKerHn85YCmCru
4tBbtUl2Rt1nsaoxIg6TfwbbOA2f3Qq7naPT1XBes05mBD/y9l4HJ5y0W2nNYDhA
WCUj2JNQi3rvVh8tGeg07VS8xXoyoma1ToOlETjD7MEdSu6S7Cw2NbUft9BdqSNB
ILb6QLTO55J10S6bs0fKKM9xYQCy2+gmY6hBKwBfouMsPqCFTupZlvVvfzYcInjj
XyEcDbxdKq00j+0PXAaZGq2h3sYGilcIZWiqEAgbn3GQIMm4UKf/yNs4TvDl89Fr
EsFkEzHjSshIcBO0NUj0IyKv8re+4+QkuaTsHr81zeq/3oggIIzG7T1lWzJk3zm5
UvuXvcdlARj9bxvIw158/QLdo/ZvMtTXAB9jAFB9ngEmdbUFavlXudbg7xslTbtr
xCjtRjiIOrd9lxn+IDmOGs/yOvQiuOcB6uIEzIWHgnF5PLf9kCI66jkYJcY9q+4O
2njE325Bv3yhLB3FCG3gdf7WevzDgKCu9FUV2uYwcX4xZjE+29f8brOC44/+Ik1J
HwFWqPRvosUpAGVhQaRqgsI0zVPfETGgcGVkqHOIGlbBy8PJLZthhneDo8oblaGU
ZtCq07+6YS9S+RvH+pZS4di9lpySIj1h5GkTcd8WkZ197ug2zEHV2OhGsuOgsg9s
Pc4MB+WsdZymJfdcDroSizJM8qlSLNDiuOa73QmZ4CZzymrjpONg6VIrCuKUPtjO
khIb620sX4IFDlG5zkdjN8k9PSEzRozu8n17bCa91MlmFfvn0LDPbGliX6sGsADC
i2O9VD9KY2cCFrhFIFNxRDLFb6Wa8yZMRi8VSLdP28GglwT14Hz9LfBaEKvZWd5g
hC9E6lbMUmFc+JP8jnj62WHbDyPTYiMH2oG30uo2/I7DskorhIp3YfbWBDd1Kn/Q
mbkcf8ONElY2C5G2uv087x6EoB5jNKR1gN+/jSSF3aWbtpMQ0rrJ373GfeZuzJtF
r6zJBR++NT3/UIZ91XFjn7ZIt8LWTm0qoPXN9i445WpSVmg+GG7tmauSJ6ebTcct
Z13XxpXPDweneSxNDwCiSWuBVUkbGQvqXXIbA+tiLMdrBzkPOIUsSYW95+hd6fQ+
3P/9DS2qdaCTRQFmGmDuow/awS5zdbAhhaZfpO/ozQ7KRMJ3VRFRfeha79XG8KGG
y5zeej51kEopoC9BPVMjyklvTaMSSmfU1zwWBwDh2DafGqf7Ifv7z0YobhPvXGOA
W4L6tUUlmb5hy4sM55setFFSEQYGxrEosqcWgo0fwbdeJVgYGJHSOuLou9qwrlqH
LLPmePbYRioiRMabMRv+I/wIioRkenpa+jqb6G7PFpYDNm+aDawN5njOZEY8MYAf
UJMYOsoUVsby2NvMqj6wu3urVMCBK1gIYM0wZBAdD9waub3SNDfLTwSy9V8AwMQk
h/JdgmA/skwvnq2754U72Meyh8aKgR7T8Jpihfh9msBub4ETMCNViddro1Hf46W0
4Gfey4YdnUf527fbNgx5tElIR0rgHSg8O2lr/ceHMCuDIhwXuHtIkYovADlrCf3S
zJpGwwfuRYI96vSbvOshi11kC43v9xunrxQK8CUb1zapYNSv7EQJVSIQfoaqRy8B
nZk2TDzycAP2mVFaipZZyaePMZpvrKWwnoum69jxeNe+eOnRqBdWv45idICT1wyf
nzCq3V/Asl+kvhust/FIoY2KgoKvPz1sj4vz+gw+JwwXTd17fNdb7cCzu9yfKBpI
t2VK+dklaY4KYGYTrHnzo8y2FItXD96ryyy9zT8sioRctNefbWnQJNIdHYask0fk
u8e6KVoHM/LWCKaJAkiAZrqlYLPflIZDj6tY5YnoSAppym3+BQxLiBv8tohYzmOT
pYfZDLFzWRdOIw/YIR5Ya4Is482TnRCH6x2tkNrtaBGzz4uN7xXRepihOTVefnsy
oJ5bxNgy3SpJ4JwiIN6hrXcS42ir4Xshh2dHx+5D+VmSH9Qt98VOHk2TqPOHANGT
X5Gr/TcbmwQ1WczHjXL8CLaEAv0LMeQ7/N0EFQcq8LeTGwuhcMRpJHGiN9zz+6U3
dVa+kLrmchvhJ25IBvPzXgXZonAs6A0M4JiyX/W212LorqGWsBVGTfLnsdZoRkjG
7QI1uU7dH4SoUgvDl8Ipn8vti/j8sEP2jeud1CSb1cJiWCHztZxGvJem/VUBeo/g
/6CH/usMSggt8CkEL/XsxG8jrUjG3LNB2lAcg5RzqGWYbsh/5vQRF90Joj4sil5e
u4kQCXQYWFGJZZn5dXZSmyTWab6OHXZSm7QgwGqLh/zjsFyTWwiT8bIjPMkBYIBi
c0bGRaESXOoT6A6AZCPIyJNmrYSjVGjRyq2Orul76vXd5YBi4eVJiDs0J+8ORfEU
Zu9rEYgKIkLgmxIciJx/1fcXGqZsv43MrsITVWHFyGBuRs2Knp+x/LnpZnRY3hPZ
aBiFY07gEA7aPYr1GfkLTubDjRA6NoOE88hEZp6hnZQK5KUfHJL35U302TJ5SzaG
z/n9dvSQ1NC/l34taoawDii9M91wToIfT7EgUUGozfbJJI/65B08vi2Xr1bPckRQ
/F+rq/EflMzuYUtVvIUN1DYAKYolFWQYwgcBjb148MU4KDn2UG7yDKvkj6Kh9Tdb
VhJFASsQWrQNCGK/RmT22DyryUFYWYWvxpC7qDfC5ja2xdpRlCXaCTFR/tvl7kaa
2IfP/JJgvi2/BUi0j3ilBW9W3M8PRwGtNTwe2/LdmyaU1TrZsxr/bUVwfPI5Oakn
0OJBI19EmUmPUX0pL7B/AaSG6ngRxye0l3xE9ueydFirOanLvl0gepKDfw7OlIqI
AuLiNj9FpswGzhPLf+yexBweS8b6TUAmCke6Odyc15tX5MIY2RkTUzqsuXaMsxlB
+mfJTWgZ+BT20VOmcjAIT5rLhZROPhj+SW7TK+Mm1IAubFrpi6depsik9zs2LpMd
lUS0FPDx1fI02qtvFnR4cSEWTJxbSPy0CCYHhJPQHmJxdKZCas2V4oErZN6puRf8
9YYV7wi3gftfc6ylqZz5VQg45QrXg8vMC1v8eK7F95kqgW2vq0bzaxXZmHPe6SHf
0sdZ+DFtXvKjQjKrY0DUC6A43eIWV7dxzusbsoKrUSDq4TqOSXvn0ChihdMm2MZB
Arv7FRBAhfbsIolDmwJm0bvXyJVyhbDCTKUI3m9iSRzqIbkVoQH3iPs0wnSqXtja
WOEgTSzThubHAIjDo5/SGpPp9dBHuZOSzyr8qvR4cIXLvsnoivgvGaakYhMEu5AZ
P2xIWUgMcMkxMOrzd6JOTmpA1bZKfVMN3XwRZ0qixLgBWGTmoTSccWSaa8m0AXz9
VS4/f3MWcFJvX64WSI8zvjVvRlA2/6GPDXHCOkoGUNyJ1ngNggiWZFe3vlabppa/
a2zhZZ9BfkylAam/YyM+2m4rflApTYYEg8S4bsv49r6bfPLTR3ZcQSeTOZBcsteD
KR5HseIht3XS4TIMIwqImzi18VviZKZqJEnJRfVxKnFrq9cdXgQAd9ks2VHrNTnk
QH4d8QDugCeYN5qIRwSgYubEi+v81LHZwOLqCJUVlotIShztTyEUSsMsyCnrcbmR
I7wG+Xj9nA4uruCJnMGREL4xB+2zHYZRPxbCpUKbAtt53pts9orOBp0UBF/1WgLJ
bXKCdIzkvDoh3j5An8YxkYh2lLhA8UU92Dd3mKCcwmslOHRHMEaht4/WVehn7Z3r
XPfFpwM3UIkfzQ1JDHfRbFaO/pkka4oQ8TH1AXs0L+sWKmWcWPoRXaqwzgz8C2WH
U9M8yeWdlJ1e20OiE/TCpceFY0qsXVDTAAcQgh4fYynvVyO0FZfeEmteY7ZRv5qm
0CbJL7tglS2KdsVrnG1Uzapj9RNqK9ZrNJbm16m1dHeGSRJWgzHHdkXldzoWIKZZ
x2bNChwKxht7T/riKbs9tH0JxrR59aYDztfZBCAdTgfO1DDiFWHSTOmgKj4GP/UH
nVPrC2ngwQ3evoc9/anJV08/mm11nQrM7UTIu0svhMUbndCpIzfeHcA7SWbH2ort
YPUKVcFJy4NYxk83SGhJcxBq5mUhfSE1zZu/4eppA4Y8gCG2+pKnj5TbygiZH6RK
8BhomFi6ZWid9QLQNJ8GcUp5Ioq1EdBn8z6ISygiysNW1cBLFyALsXTS1wJYKYDk
WTKCZTjxLUfHogFvhvo3CED8cQJbB/k8c/L24/y6adoran3b0p8pxVTwR8DEFGQ5
bIM8mSPZEWqunOKbUU7QJVcYuJAhrhFwWqfRJuoTV1WLEAwtsjpeVGH7Is7Tx/at
hwyTLWgUGRm3zZH9yPktHrArKbwGllZzkwrh7VvvH92S9aMoIC3CcxrQgrEBGWZz
xGXT17duFreGU1Xuy+h0lpSuvZuesnYjEhUfTVF5G9czIMh8m2AFrEG7mYLFOKYD
4ZIxn08XxHU9NG+ST3JLKN2vfYo9/J7HQaPI36h26pgQhJ0/gL/Otb8lLnN9Dlfv
Y81rDW9cs9dMNuzCbYOtsP51UevdJM43uqkL1rXWfN+lkY79vSt+hBTwK7ro020e
HpcxOjsQFWF6Qtn0vMFX/6lp7R/exwinfiKE27/kOUetzMkvDRZ+gU+pSJNXkXdl
Tzoe6vLaq0v5eDPlEcBGXz9GDwi/qVf9I3HGU4XrNc6fgXtq2E5ZYa/9prYJQZha
hgrFx1i9wRTlEVFkuAZ93uj2DjjogGjhUozuAjAdFa5f+cNLA8e4Hozd6Gf6Nzba
VOfo7pV7eE2yojEpdY9s2cc/qK7Jp9UL0pq3KnAg6EiFoP2B4VL/n5zNnoJO8YxK
w+fHSeqit5hXNihXQCMs28ojdfxS+cidYXO9jmowTHFcrrPOJ6+OmIB8kQRCMayB
XvB8XDiCccA3xvXJqV+mw777Qj1pC5emtuJXKlJuTdBJ+i+IfEPsqvrTuQznpQIw
gDahKOtPDznxe9U4hAnVmyeV+xHo8JIvtDKXhhZUjYB2dg7juwBH2JWBOGft+WIw
dFFpG6o5aNDBZ70t74erkznXvxpnav/2RfDp/gzrO6dgaimsiBS4Ab7dcSp4+9RX
Wme+z+0eFsq8kUQ5Pscoo+g/yzEyqa3vZCAqS1tgRlAYsOf69qvrnYvoHbLFvCHF
9Xr3d4T91KsTzZEhihFeGDmx7Pgda9wveEBNttOoGtloJRaUnr12IhToUyka7mjt
SiT2xmZdxnR5t4dGI67p35oEk8vtFL+ggrRZWBsBCdB+glXDDvzg9adz5CvM92++
r37PGhTbezfPyLPaLdlXfLOSSPwPYZI8nJrKFJMX7sk8BANjuQHKmRnTy2QUH+SP
PDybQQJEwzW+lylab6slDORud5C5unu992bPgaXuXfciOytzfJaLt5FHVqk3ivbh
RzmRmhhq1q/KqPk6wwQcVVtBs/rDrB5RZ70+cNmCH2FHAoCoWlrPJNrPFJTGcsNz
7Op45+PxPpz/JRmfBOXIqSigg2wc7LYJ9r0tyjctH05Ac4KsehR/XJK95ZOcLzbc
7iqYaN/b58JewzqO35JKIPy0VsM/bq8Ds7GkCnx2Oph0+67CkcL4XHTbIQxgtLih
ntHuA1orFyIjALB8yy1jVqoCtdvvZ2xKC5yzHXGsT3Um2HokK2x/2IRQ+WcwP3M+
Ez1jPtiOMh1B8UvbHw9s1mcRmx5cIp0wk84Ktr8s34LvYXEbTsuz5DuG3Tr7Lto9
wtLH8uwr53aPxMgxJLjwrDTAFGFAHVLRtI5KN1DS+Y1l5Oz8pDv7EZAy+MWc2QTZ
4jbxcfZh5QR2msQ/LDYlDi1IoKD8tignJaLK+UQNobuEO1/9yM69eYP8zUcCM794
aWh1qT593CfxCvR0ycJg+8a/J6YfWuL9z5FzqeQ+dxijpAVbr5WilssOJl1lh4zr
77jL1ug2UsIC3Nv/zLyXzRBtdcQiK/kF06dMD4iDnJFfAjf/ZCawlCfO8yqne187
sitBU48JqCHIP7pEkcIDhnJ9pvui5rpT13VNannjiZ9FaoDkKo5J31RWCP3YulA4
xwl7aWzTn51VvjEaBQ9jKdxBMnKdTQQGomn/fcEe/YgcY27dmraBE0lmvot1WftZ
WeKaqn0cahIp3u0dE3GjffGBOkJF94zfXfy0TK607J51IyJKAmu285uFqChQUGeD
aZQeAA5NahtLUwUUKL32fmdAYG27kDA8LWa6x0mO7/UWMRNhr6QCIXu6yQbof4fY
gonWu1Kc1+gor/towJ5qdKxjE20jr/ERFM2sGUr07bsdy0st/zVtugeM5PHnR8b4
J3Y1fIqdb2Gtz5FMUfOlo8HAOETl3E5Axxqp85h5s5TVEmQLFb8OS0gA0qOak4+V
Y3C/u1MS4u2z2MjHG6MX7DXDsNaUpdpKcSXJJTxXw6/yOsIp430H92mG25c14KWF
JAhads0iff5XWlIxcUoU1sah5BG8S7gNsAKa0Z4Rq50awmciaRRhAiuovNaK778e
PaIlgjJUukuiRJsQ9sgpmAbjUVLB1fLY9AQkbgRORT02y7HZ2LxrtLIxyYjACHD0
HtA/LUr+/P3SUpEeHsGtP1oDB8pgn2G/rmxKRfv/H1KAAdPWj6vpUNiUbF6dr2oj
IY5Z+Ju4pCBNrNNHz8ric7Lc9YpbOmIP4RJIjq+1FDjKUqvHEs6aO9LiD1R1jcom
B9cINiloXwlS+2oy7XnY+3Uv7KljGpYDhk4V8wUWNwb2hWEzAx2hBwYgHy3pA3si
JR7hdj7i21dou73THrHNGXqNpcaEsYC+flPYPrDT5K1Dh1pkQ2ip8r21l7JU6FFh
9YF5AXa3Oq/c2J7FppVH5h51mwaJfwG3tybDbF2ZoXbwgzyJc5OTdDEZVxSO26z9
J62IFu3BiJF2T3AfnktHK0lVVQv5tMYnkKHqjw1sfpTH3ewh95PcrTdBFxkJK/iZ
Lt7yOJfgklJUqnw7yxkoijUEOJJbeN9989XgducMy9nhm4K8Hfj1E9wBW7GIIPvf
Z9nph3uGgvDkUC3nsXZTAK9pJ89cfVoQl5/Gj1HEHxJnDeYpOWNTMy7RreRMI/tW
uKP19nNhfmmqS/ybtPI40J3lWa1glvDHJFvv9lzVBCVO0QOqoleeLOrmv9bvFO1j
4iDjNFDkSMFmPVTv0yusW18miE5V/Nc3fO1YKtz1MIpeWhRm70ldOH1fhFDzOcYu
+Iv+XmE9cRakYEoSszmWQDOaHV6S2vk+ABlLo87zNC4gSlhvYcahr9ag7lXOMlrN
1aqUWzyMTqCUCMTg3IOzKvvAdAQm+nkpuuhi/NJwEmgVFLYoFiEIkzV+qf6H6kyq
tl35BIaHW1fvZy1lLQEkB0HCUInb69TOiIqhOsMd9pe2y8m2taMXAWxOReAe+IhU
Nkyh3IPcx5ezbhqXmnXcx++UZieCZ5OrP78Z95Jv/XJpDRn/kMEW210LPC6H5jP0
Hb5BBL4zTcrgL4Ja37vwtcUr7fBjz33TYKtdhMT68UGa4+3/rLjUzWpAeH0dpY0N
DU1zZsQcq2bPQOlaANEhSwMXDOKoeFQU1VK/tzo/HsEhI8qAJZh4ZxgjzrA1Bqgp
n9MDWFTBmwQZllkFl89zRBSAz2nCPQd/0A91oLO4yJD9IKQVFjDKrJ63M6iUU0Ca
jpO72+9i4r1aqZAvb22iwpmftmlbHaLP7wc9rmcDz9Poj5dPDdzzuowNkeyEDeGV
UHBX3vl/iECQbHRlhZoCjrES/SX3axkRnO4EXhCduI4kJkLRFJ1d0VWozbUuU15E
DrppgMTep1Uvv083lyShb37BhKLQJqgWY96aigRG9jYULMzWj4xW/sIKYHoceAs2
54CvK8tPCiUkMB+3+sAT8BCK7k1lGPGL0mXzORVCDrKT7j2p/X6EyqZ3sCZCFqSb
qn+nbJpnrgqQy+Z6YyvebjRxmpcpwEUQq2+LCp6rY1E15Oifng7SrMPhywJNBzIP
amsZHpMRWXTCdCFkKBZsHtn5nOQKgGv2Rfmxynqdpj9QeHlB48uiurxUHNwLCydz
bIb6kak47dZwuLiBZz3Jue8fF6WXsPYw3F6VC4nQipYe8d28XpQQ5Fp8jSIfm3Ta
YYxM468btlDwJzhVoLZ7H+lzHuGBAilXwPunPcbX4lENWssanrfiD6gGyu/1y/pt
XLaEKlrBgwjGmqvoKOJxHxt31Eyu/mIyknFwWGebWc4OcyjSVMQEWGOlxi9AhxB7
WiMbDX4BJaZ5iU7wlCCxgSG6y9tIGJx0WASK5hqR8s7lMD3haSJb9md3dlDD9Kke
+c7x4ziVf/CcHzH2XyfVqUd7Iz3ZZQ/W5XmZmtncNfrrLn0XY+kqykkN8x553V7n
Cpmr8gYH1ff/qY+ZVnmrvyJQfPimnqQfkDnlRSFuuj7g/v2TszW+NZ9j93l433rX
3jdBDO5PX/ghcJeGHUikSW4GoEGipe9wmOwjHvd+6RnylnXYJ3wXFN0hi9i85ZC0
8vWgq7hLHulkz8OtUkc6uuB/OMPSVneuPcSehLoaaIiQKb7HY/apt62Nh6b2YmLa
Tsu/5TSjJJNtgOYBVGk0GixQMTx+C87uoNoVdmC4rAXtVXS+dL1NGRk4WTU7z8aT
7qSj0WHh0k4Q7LFkKrsynQsLFNrwYAXmYy/ArThvRcI0ivDnOoiCBOymj5VX9CJ4
G/A4ZQPOr6+rzF1ZKxVu1aTeYlSSznr4eg4SzHADpOwMlKsjKDIrZJInbZEuCV9R
ffd4fX3AotBAtKslk8X2afjL7+78ALAQKvfn/N/0MhFNJcMRYrliRy51y9nQsIxP
xjJbRMDRk+z6EPSqe2OTKyu67PvHrVhk3mLj+f9p4cVPsd1p3Q4u4L0dikrUqLjw
FTmk3wwEuXVjWhvlPtscewVA+y2SgAAunRSS5vbrkM417NFCe45zFCWr9ANUICHn
u+vkc6PjGp+2lBPLXDNx7jUo+OdEVO14W9daJSiDXA6Iu/Ph3KI5lvMaPCRoMW/m
Zy6gsykyvDMIU+oa/+SEgDH9ilkgRMZO38PUVECu/VVXmT0g9BJIBTLg3YC40Bfd
0NnPG7IghweF3RfAqU5T1svwqvdVxT9O7x7IRepsRJUD0RGoZp7JVX/Tj6yNyny8
b6NX+cLCmPiJrWFQAPVQPsdhDIlLzKH5SAO4fKRkvOB0acz3Cj/je5d+wMneQQwD
B4pwsNmckjKUVqDeOjiZeFtvlTgB4YYN6ReeBu+dWpq8IeOiVQF2wzGADi4sbrYn
yjEaIDkxyucKbELaFH/DkzivtKh4oW4naavSstEsyrWzotzvFlXYXYAOct+iSjyj
N9sDjBv3f6O8rq3H5+5larBfGS9FPvM958IEUYMGoUQMGdQt9gj+ohUsN7EB53ln
LBzUtzfcoBS19QMHO3L4zUDT8COb0z/rtYxEN9Cayj97fwZuvPgVgGEIMRjaeqLp
NCcdru8vRNDNYvRneLi2lnmBSnf/T8ycPUqqCr6lqlmbOUFeFiMcgAOUP5joZIqn
1BIn4+y+VMBDlP6fxyQKzrfGbNmeI6V/HaiUURRdHGJhKdpm68B+nxRYa4x3B/N9
BCv5fGpITiri6xFDdGIAMQNcxL+fEAJknDHC7WnZd/whiGmIho+7UvXfFNqqgEWX
vBW0xfG3+Amgd51y/n8UCJgmfStCZrlrmadgxfQRkaaasRW84A24uIsR51ImzDtq
9fQx3+VjcBDKnDSrOOrgH0JJBwLikHy/f52lMxT54pyM/QcvWMBryaRQHOCjvzME
oHOPd344JCLmIN2Xp0EuKMeACJWQKjUjfICbnGLSvWPIcUS2798yRlTDv20zabwt
mxOUqiMRplRSu6Ym6rWhPdtwbhvMwCoqYTINJASaJMf8CPXni1ICoABdZs7sBtGa
s7nVDzMzU6/JFcXjwMbohpMr9NBpVtQ/0XM9J1JWvx8RgVYKuS+6HJKhI01wvneu
TRXl6W0cIfHTRRzfnYugH3uFe6m/VxKLsvCVmqyL07DhfTbp3LhLlZydAswJ6hfM
9Mfh+u+5uQpk/u55PBD2NcMaft8jqUZxPFxCfiKUYy9Eu+TU5bH2U/x7+tB2XFha
L+5UEOkL/Z2vVx+5kJH+EQGXRgZxAGVdqaSd2jzJuE9rrCbSk2HdcBd1ZwtxMM15
HpzCcx8SH4W6spx7iyT0OA3K1RiSlmcAZ4tXWUjgC4kiv5sChIjGnzBErsjh1Div
GAgBxoBsVhRrSYbLmXwqbUBO4a+bhH4/vOmIcRXlkZKoKl8tPssJLARp5sQwOmLD
AJkqxBWh5sI+v6YeC5TKJUpPMzKaAQZLN4ipUnO4753YkIa3omXZHrQd6biiFVD1
tr5u+imFZeZhpXfPEBbsl1ixI6xtywnRdTgyWYOww2Ukih25vQ13T9xVeRpOzZ4Y
Ew0nRZwBoT+q8hbmh/3MH2UNxxdz8uyb9EjdlxNEK96XXGrVbukZCvCLCOPyFJ2z
NYNCYyb/+iADnnWf4XtpwThBeChyH27rbSTA83cn5jjq4S5YGICM4ofwSTxJOcuF
LIySaYnfPBmP0rnArJqzIaYXY1NzQOX0F6jnZe9+waCjlv6yZ8z5rHnqpWmOQD8E
nrEt3kzWP1dxZwuzaBuvXPcqF1Ke9sOZ1MSdvZnS/qnNiVTr7Nqyu0prOVUoctZv
XglZCdfK3MCtkEUHYPpOUHzcBKTTSWrj2mzbGttIxppAgLPdJDhCaWmJbB0v7vqk
ytcDMW+5RJ2i3FVajZ/HGXMEIbsfuounr85t1XdGw3S28T8S7D+BK1mee5MDBV0J
lBuX/Evi6JFc31luv3kVAkCQHDkBC1aQ2Ih/QX3fwAoVw44nI6IiwkDaVS2gO5Bk
p9qxNB5JpQdj1KZJQu1uB5D1DyS1DDomLrJIokFikzsuWun1QZiEw+CN5xP6qKFv
u7VdYaOCNMG3YpzHqs0z3/zS4C/KAe+dgUQG3pc4ROdW7eqolsvb5u8mFeLfIKpm
lMU7597mrSLywca7B4xIc/ijl7npmg4oyx4Xt54N194pg+CCFbXIMUNS3Fnso/EA
9x0pa/1PCu7GB/RxfxB6YuAwbmx91jJXw2XRAbj99GQ033Sm/E3NJ0+3fAruYdj0
gu2MfwV2vUoO370gr7LqK3c0souJ7rJR3CmNwwYCx79lkLJztJNVrXDvSGS2rcuC
KqRpYpNkicf5jPdjkt5plfxBIN/V+Pd8FZ+l/CPB+Lk3eruh1C3P3ZZ6zu9oZ144
eYi9mohnDL0KkG4lPAjk03jxN3dbr9dSXbm4vc77dLVu0ZC3rgYRczQ1DrHMKiHB
P14drxKKknnJjjAx4hzNmY376PflP1ZU7oLliDmdsLCu43YmMs23DR8VE533QbqE
kK9+YMNDzHkEpUi29o+ukuk5u/K26lQH9YFi7o3jYnQhazlP1lS1YvpoR0PGa3xn
eQnQWM9j1dnW2/ElR0LuCa/a6ntkcIjd+1UMOopVSvllun9liGifSMMF7aiiB9Md
mW9NM2YFGoFi2RAoqoWtf8cULlzhWhTdOrOwnGfhdwf0J0hCIKQI7Sjx+Yt2TBIj
vSDlM+DAgzkDVAlHwzFZ0Oj6tJML3YFhFmTTB8CPrETjr0RUTRO27dgc6pMjS8X4
XDG8RcKtJyFNDL+qFWJ8apqIO3vJmKp+4kXpZoCUqS46xtING7xrWL1fDaEMAc/F
/orsO0DOdlhQilN1u08vq1t0NyhKpstzNfCPjQTvc1R1YLnMSxXnGZ6AwHBwQ8RF
Ts5qutFChPY1F9/4tZCSEjhL23fLprE4fnfZFCudtHWveNHpEDXIlRHUbSSFtAgp
OkRvVhhAxNv6WqINuJEqq3DhyNAp1UByL8sRt8cqIrJrmSox+kV7ojXABeMWi+g0
LcnhiBElAwWDW7sV4HxLpF50LYkAR4IBBJ8HRzLN71A/OwgZQjMtm2AxMqJEr7l4
I2EN41HPyto4w5Y5DU9AndWuizrGORbJ8L2TX2tpQqzgam/eboY2Qevm4eLwAggH
RApODA+hnZiaH50Gb9YpeqRWJg2DFwEzLNSIcG95d9eO5AG1puSllE+Ci7JUToOI
/H1/9OWj32kVEpuywOSJYWQM09l1h7Ryr112IeRVUqcQgZWnmc97en4zM9tFte2d
7JcmUy9TRiIcVfW0VVmc3f9x0WEtP2VuQCh7tHM/OuUW2EAVZ4vjv25G1h84kXTS
Ut5YsWWVrI5/tQlM0GrH2BCrOceQHR2rqYD1gpuDakkM/698aTpZy7eNxHLHlX1Y
9GpeblSjK8VLZBq4ELszqmA1JSKToIhrBkYI1Tt5f3RJQJdZNuco3Cn/doCNn+7I
wGZq+oRrJ3nBuqHKozYZPTohsEmf/9fI57Ti9Cpcj+4M8v6zI8gXY+MrKLUIEfOu
njRFiuoaZfHZFMjRrE2jDN3BYCnBLc+qr0r6iyrrcEJLz31Y186Myn8aMaE9JCo9
QWYbUyBiKwMR71ELdyxp2zCy/mxHnM6PBkZZfCYfs6c86hwld63Csr9sl1AKprQw
i9rInnf4QeW5e9+FKyA3NBoOH2FzuYT+T5oDP/7lMOJG+rYf8dvtm002aTevBP5V
hNjWC+cjqazL9L23HyIatkgQK/cfJc0iWf1lZIwOIdA9B2T/5pX8mQyRDRSLUXJn
lLYhLHkvsAjJps8vlv9F8+Y4Kvs85I5FfCaIlItkevd9Lm7FRtTjQ3lXy7d4QTWW
ekhtM2H7lGNn5a0NUugwTpvPzkOBpXuYLM4odIcYiKBgVN8dUkMRnp6VmkKFnPlo
zJmMHkqizK6017gdsMo+wMvhNldOOdp8tax4KX54ZgMxEBV0wpkzEHAw12xjvYV5
4VLZqXbnRK4WSBAneHenPYCN3eivmHMi87VVQmBr1xvJGahP5+Z4TpNDSA3agC9a
D/dENqV2LW8MJ3mnXFvPFRvuewLrwJfkeNREq9BYuepceXEJ+nCO0kfBnauHF4+9
c0DgODsyO9ChKLuk0RtSTubUOlYeYp2X7sHFXMphEDgvpHAYIfjNBLEafKSaZvrP
/hxV8LgiubAD09YGE8fGnej/z7qRC3+1t5SKLVB797PzHdBn2kzxsL4dqNvT7BSU
zKQFCHgxVhsnUqp4u578eah/zqZW8Nl0lEHTcbSHaKYeyghluuNQVtER/WztlrLq
7GnNU/knUV8K0NKyRmQ7CZdgGefXWSjbA09QNN6PcDNbsKOtr47DrANE/Eq42Dgc
5DTp/8zuNx/w+/qd9r5czWeXi1uWunFN0ZhL6paX/hPBWKjNVyWIDveswFjuE9nK
dJOk1FITLjT/GPvl4YD7Okth2w10GFLgUMINFAE9dEejNh47xw0Fp1xpYohh1ozH
w+mMAS8sYN/fz9bf3cYK6sHe3SuArUOqUF6tGQ4LfeMmiXqmGb95VcyE15kM9i9I
hAsXH5WWLDaiHE+lAtxdpUbZYASKBmhYrSD5yN8nAysnp4MHev9J5JfMx48rFvRW
YHPO6LIhqTNfmhoXnvutdOxidTQljvbBgCYJfu5GVjFTxuLCdPzntI0B8RrFXp9j
MinfHGkfq3eEShxMcbDRGoVEjdR332OjGdU5pw9Q3UjfBK1jiDOA8XeqA5QKZTjr
W4omYD/8EjjX11Q/OXpYjIE+7hXeNfA7/ZBaLcVuI88szVJzH45+5PyoHSYdNWeA
/KoGOJcwxM18EbSup0JPV9FlqiYwhB7esK46Fw1MlGYF7SDKreZ3t4JekjvIUWxn
bsDdWmgqJclDPZwnTJOB/9iEA/RHCSXdMSDEagFfkXXyCqCo0bU7ia8vs9U7uNvy
tu3nN7Rje5A5x1z46Fs/yyv/DXJljqf1W9GaHp/b1Gr8QA9wjLFRj2aXDd02m7Yx
I49o7DCV6OCA+6qrkDmjCNQfo0USORg8hVdHFHREzv2aJp20pD5EdZ1Fudp6mN2r
OtCUShLFGx8DHlpqkd+6ObVd7jW3jljBSwvQVryO5J8y7TCxH2qHcj2YXm5CR85F
t+WxjxAlVp2lCVCp4GuWpA1B11g7gl5mSYkbOOOSbD8imtTPkL3f8cdxB5CqUMYQ
Uyoivpo+EiEeHnaPPFbbumTUdMe32hjUVTasjv2K8pfZDYqkmNYHG5AgZYQKUGSy
oD/oDBY8USAmmO6vD6H7MwO925F3v9nt+0x8v9WpPG0pFnPdam6DpnnI5ZI1XHXd
XAx0jAX0+hAM4dtfWfJj6fCaek/vkIh2yTq8KYypKriOOggeOxi0SsZMmvmwS4SA
rU0bR+BVvWMdIaIU6541Gyt75AG8RXO+gqk9yBqWYeAv+NJYHyW0of7PLBXCsNgu
w8AJJnnZuaC0/ud03TbN7XqGO2bvAVH5fh68Gdp58/1Qt5959aFzaNB8s2eyI2JS
WoUqQ487HqfJR15zV9Lt4ZWVxpFm+jFHHqyEMk6ZF8IHif9mMCiovbd25L9mxHxm
y/tqmOQWvMYF8ovM02SjnVHjsd92ZauWRxkCjc8QoUkVqCGjKoVm+MVHDGjdEizF
TGy4ZpCUsy/N4/3/w4G1mt0xL5MZ2/w83J1SVPMosTRrdelPovKEWRYB5Tm0wG5e
cK2fPHnPQ0r+7N2ckGduVoGknRXVEsEO3Hz9n8ic1xerwOv4uaboAKN1TMwROrxL
nl8jc1ALtxlKlEk3kbXj1ecr0m00TXnG/9m6WkuBCyhDbCMiTPhbXVrFt27IjnB1
PraRP9RWE9RA7p4NPx8NS3TUZ0KL/tUYbToKG0nA2GQhUAWf3osl/GIIWuyOQ0QW
liiOa1FFQCvmjRMnL5PIcv+c3yF2DhvAaW88/s5u3rIKeua90u55gZP3dmV2ixXP
avuUuWyrEKok5fOWpB4xm8HXTw5oPxGUVE2PLX9qQxlBPFnjSn6HWa7HzkOJUa4a
Fcnblcb/+qGXCc/MphmQowdY9HwB/YVpuXpN2fdxZNvrYmUBSelhMExgfpzxOnZE
n2lWyYrdER/6ibMLXOuoyBL2H9launCGioJ5Z8IEmz9PhiJNPBtfYU6lWQ4bej5d
ifz1+Ou3qUo5CiIZh4/I5LaH1xqBxLk6o+5HXEWrZ5BjIF/badPPjhr0ZPT6NV5E
M6K/zK47hNxKAmhnIevxmUAbsroiRUW+8GL+rBqIOUYEyd/OX83gsh8lTxPYK9u6
I+i4S42ZeHp269fR2yJPphULqRaIlLeP06ticdw/E7Fwja3HtgyVZSBKCzqdwv6Z
+YpmaDyOg0imeuEUR40BYun+116ndG8z1yenPXCYy3RPFKrsjEA+RiJ0igSVGr1F
8mqkWWOo9/2uYvW57HOrEkRXXLj1qU94gQAS/4dyPtJsNBPjLj/YfMB3fmHCWQts
xrdENZ8Lu5mkVNJc/xmFmnVpObH1UBD4XB/1jIa0gk5Ij0vG9SjGw968YsoEJvtA
/v7oqnZwgOmpeME7ZMF8pn7mgaxZ4uSIUl+aHg3gUAzwkWv9dk8g7TFDhObi2IPY
vdeSHCsq2y9aCJHvQuzZ4z/c5HuDPOitpBJlhgbYzRKjSneDkxE/owXw9MaT3rKO
XUYmtAhSCpCScHAsDVEMc3JynzI2i0r7ZtdyjSlJjvNNRItrNOkONKDbQHV0mBj6
UqBL/MH6zsD6kwNwlBC8i4PvWZ2kOE4PY4/GKMavZGEjUiH3MLlx3RLay+DHaWv7
bZPfflxIuzNUtyuZ7Fq2EvBJ15oZOnOqdztw3teKBw5tT7IY1oWJH3SAfyMJ5M3c
ky0sYtlb1qcUN18nKJ3CWPJrEwnGI4Egm1pqCMmkqh+Of89aXh3HTI/YsGza8iNA
h6VO0tIfIzRsQJXXaXBCT5I1KumNuwOThNoCd9U6WUE2OYf0ENLwlFAQkgBFH4Je
MQjlf7W5TUXa1bDxlGzo9pnaHSXk/5d+uumsi28ywEFctop/rA1vFGtwiY6idSuh
eNef3gXZgFmwMVOciJGH26lv/+tohNO4A866zMnOqWK9aQ+Q3s+G75zmoSKBBQUn
QIzf5tws0FeYdf7KGybH4Ud7gEjIo6dDHf90aR/FMfz2td/3ZXq70we76i6NKWcy
946fRucDUq+ZMEhowQDXOEMTvJPDTZHba7MIQwgCnELy7YgusqSSpQlBhXB6HWmb
q+qmHKkan6WFrkqvTzOPRUJ/7RASaqH5JIPAxVzIyhFKG0E7iHsP4Bdw+1Pgt3oR
mCiN9DirsMpS7ZQ2aZvl3wmy0JffVI5wP6kaJBsGC5xrJaNOvsmLwjI9LOEof6ZR
UE5iOrUbLtfBBWjhL9EmUoA9UcW7P0f1qV6bABS4IU08jfhCiuIN34c2oqS3WZcI
2cf14AM3Lc+waLF1HbSWocaDlaLJ7LjDTCqQplatoXmFrbvKucyYoMxrFeD02AKz
h0cffaAH2PLRpGq70TheV4pa17/7qDfKCgXmH80F/3Xovb5PKTmAJgeiYAVZU20P
DUKiXsWVHBRMhm0zTWlX8/QS3LOUf3PvBTYrAIoaoDhSa70co90Fo33KZ2oZWkxp
9VEgxywYyhYf7wDwkSvjRj/qMv9o7HmCagCE/U0h5wEv7m8PFU/Drx7Ionj7SNw5
wPNtC8bsPpac47s3FSFUQiySkonZybjtjwO35MeyiZnU82M0f77Ra7+4Zwo84dwB
vBftfwOSArhEUbpvSuDdfFqPqp+dr8z1owVa7+Gr55uJSADPXWc/pcArJETdjTAZ
V+dSnv2t6SgeTzGZ3ndZ48Yph9PBxwTNomuSYdoKTZ+i6Zr66ftuNw2SfegjPVzA
4lNeMfOR+lroxcvMVN4sSmGF2ggtgH5CRySjQbYnQXtiJpZ4sBZX3+4ZqhDX2X2R
Pt0LnMRjgpNxKEk9oCtT6ROXPD4d9QoyrSdlPJVHRNBUhzI1MnG4OhFdcGPNBjng
AlO3OLBmIMRRL3q+F0Byo4+ue+vFv4WsGtTLQYARmj4EqfojLp4b+cZbvdX4nbey
g6PZQNLhCRF0wMD9vBZLxQldhrf5D7j5lPy8asF+2L56XvVxiwzxl6TrO8TeRo+9
tMwc83StCwjcVLTj5f1fbjAzCuB7Y3MCSt+lHZfJpks4FeDars2bzH08SMJ2WW2V
RdCuotF+GjNHG0tQoGknnoddDUhHRPxfvx+nBmf0LSijzmhIg1F9291+cqq9pf5x
jSbT0HHUS5MvBqDmhlunUsgp4QAxnqX9xqRuwI2jFHJ9mWBMpwB/q5xk78YCdz5U
zxOAtGxTjuhqkLq3Av1sBxNqHR5rf5ExIlOmeC5MiNQQfgxXsLCbYHRDvTLi9xJ4
lKeWdTnZmQiLfsIIxZlCIuHgK2kfSc6ioOnpQSoxY7Bse6PvTyutWZbraD1/n4Yq
ORToy6P0zRT8kaTtKkRyFokU/pibt9oKk1RXct6UkhfNe+Jz0yWdLygh0XsYDogq
AE7lO1VsBb+NjbEI7K+6+HU4BOH3tJNplRjCfnDViQeWlAb9eLYREjJg90niY3tB
zHQ3UHrrJwtYinqPL2icEJVsDfV1IHt2WHwFqNQlg1CqVFOF6/maKym87XAnDYXD
DCegB6yFLGtDNuKQoWZEYmFXszURYZSezAmjvGetW6pLqUGI3Egp/U+PVjo6GE+h
i3dFF84atu7h0metKlZpIB0mPR+AFlc6t9smr11AAblPDxMbYtI/dSZN0NwEl0NF
kMqt2lBYEfFUsl763esJ8qB+Q3gDgYBsxeEDY85COMI7qkbp8S9gXq46sWJnBLiK
8Yh8GE4jmklgd4suQXrCicu8j8jKkAHk1CyUeBIUsIT8OTogITLNgfrw7WW438Ly
jHITLyaY5emQhMtjpnUqbTZ/Wgh8CaCC1bH4MrJnjIdfg8X+9L6rYPDg3cjHZv3z
P4+CIPib3fVIjvnst5zwwpR8ssQwV+o/7It3kyx6/UBRH3AiR9FLNEB1LOdJfffZ
iNfxYqZ0c8oUzZU6tpmRTHASen0l5i6K6oavTo583LoDF1iIAxLHRiQrmwuDEZWx
uc7RUtMOF1ZxIUE8CKO4PbToHJAVjnUIpQKyvKQchs2EHwY2Eot5voNczpPYcJ27
wqhN9orM964NlmrZ2O7/c/drOFo9tip0XlUN2+Lo9vGcTjMiKFby/vlKUuyCGPRK
yuED0qkJdoCQ9kWUCz4/+gQpfLlHOruQj6FTJW1OZvBK49xuANk3dmIeQms5B6So
QgIcbm/BUddmFzWk+pXh1iUElgE9gzkvpWa92srzTJs=
`pragma protect end_protected
