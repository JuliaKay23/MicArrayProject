// nios_system.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        clk_clk,                             //                             clk.clk
		input  wire        ext_irq_adapter_new_signal,          //                 ext_irq_adapter.new_signal
		input  wire [9:0]  ram_block_s2_address,                //                    ram_block_s2.address
		input  wire        ram_block_s2_chipselect,             //                                .chipselect
		input  wire        ram_block_s2_clken,                  //                                .clken
		input  wire        ram_block_s2_write,                  //                                .write
		output wire [31:0] ram_block_s2_readdata,               //                                .readdata
		input  wire [31:0] ram_block_s2_writedata,              //                                .writedata
		input  wire [3:0]  ram_block_s2_byteenable,             //                                .byteenable
		input  wire        reset_reset_n,                       //                           reset.reset_n
		output wire        tse_mac_mdio_connection_mdc,         //         tse_mac_mdio_connection.mdc
		input  wire        tse_mac_mdio_connection_mdio_in,     //                                .mdio_in
		output wire        tse_mac_mdio_connection_mdio_out,    //                                .mdio_out
		output wire        tse_mac_mdio_connection_mdio_oen,    //                                .mdio_oen
		input  wire [3:0]  tse_mac_rgmii_connection_rgmii_in,   //        tse_mac_rgmii_connection.rgmii_in
		output wire [3:0]  tse_mac_rgmii_connection_rgmii_out,  //                                .rgmii_out
		input  wire        tse_mac_rgmii_connection_rx_control, //                                .rx_control
		output wire        tse_mac_rgmii_connection_tx_control, //                                .tx_control
		input  wire        tse_mac_status_connection_set_10,    //       tse_mac_status_connection.set_10
		input  wire        tse_mac_status_connection_set_1000,  //                                .set_1000
		output wire        tse_mac_status_connection_eth_mode,  //                                .eth_mode
		output wire        tse_mac_status_connection_ena_10,    //                                .ena_10
		input  wire        tse_pcs_mac_rx_clock_connection_clk, // tse_pcs_mac_rx_clock_connection.clk
		input  wire        tse_pcs_mac_tx_clock_connection_clk  // tse_pcs_mac_tx_clock_connection.clk
	);

	wire         sgdma_tx_out_valid;                                         // sgdma_tx:out_valid -> tse:ff_tx_wren
	wire  [31:0] sgdma_tx_out_data;                                          // sgdma_tx:out_data -> tse:ff_tx_data
	wire         sgdma_tx_out_ready;                                         // tse:ff_tx_rdy -> sgdma_tx:out_ready
	wire         sgdma_tx_out_startofpacket;                                 // sgdma_tx:out_startofpacket -> tse:ff_tx_sop
	wire         sgdma_tx_out_endofpacket;                                   // sgdma_tx:out_endofpacket -> tse:ff_tx_eop
	wire         sgdma_tx_out_error;                                         // sgdma_tx:out_error -> tse:ff_tx_err
	wire   [1:0] sgdma_tx_out_empty;                                         // sgdma_tx:out_empty -> tse:ff_tx_mod
	wire  [31:0] nios2_gen2_0_data_master_readdata;                          // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                       // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                       // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [20:0] nios2_gen2_0_data_master_address;                           // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                        // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                              // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                             // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                         // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] sgdma_tx_m_read_readdata;                                   // mm_interconnect_0:sgdma_tx_m_read_readdata -> sgdma_tx:m_read_readdata
	wire         sgdma_tx_m_read_waitrequest;                                // mm_interconnect_0:sgdma_tx_m_read_waitrequest -> sgdma_tx:m_read_waitrequest
	wire  [31:0] sgdma_tx_m_read_address;                                    // sgdma_tx:m_read_address -> mm_interconnect_0:sgdma_tx_m_read_address
	wire         sgdma_tx_m_read_read;                                       // sgdma_tx:m_read_read -> mm_interconnect_0:sgdma_tx_m_read_read
	wire         sgdma_tx_m_read_readdatavalid;                              // mm_interconnect_0:sgdma_tx_m_read_readdatavalid -> sgdma_tx:m_read_readdatavalid
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [20:0] nios2_gen2_0_instruction_master_address;                    // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                       // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         sgdma_rx_m_write_waitrequest;                               // mm_interconnect_0:sgdma_rx_m_write_waitrequest -> sgdma_rx:m_write_waitrequest
	wire  [31:0] sgdma_rx_m_write_address;                                   // sgdma_rx:m_write_address -> mm_interconnect_0:sgdma_rx_m_write_address
	wire   [3:0] sgdma_rx_m_write_byteenable;                                // sgdma_rx:m_write_byteenable -> mm_interconnect_0:sgdma_rx_m_write_byteenable
	wire         sgdma_rx_m_write_write;                                     // sgdma_rx:m_write_write -> mm_interconnect_0:sgdma_rx_m_write_write
	wire  [31:0] sgdma_rx_m_write_writedata;                                 // sgdma_rx:m_write_writedata -> mm_interconnect_0:sgdma_rx_m_write_writedata
	wire  [31:0] sgdma_rx_descriptor_read_readdata;                          // mm_interconnect_0:sgdma_rx_descriptor_read_readdata -> sgdma_rx:descriptor_read_readdata
	wire         sgdma_rx_descriptor_read_waitrequest;                       // mm_interconnect_0:sgdma_rx_descriptor_read_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	wire  [31:0] sgdma_rx_descriptor_read_address;                           // sgdma_rx:descriptor_read_address -> mm_interconnect_0:sgdma_rx_descriptor_read_address
	wire         sgdma_rx_descriptor_read_read;                              // sgdma_rx:descriptor_read_read -> mm_interconnect_0:sgdma_rx_descriptor_read_read
	wire         sgdma_rx_descriptor_read_readdatavalid;                     // mm_interconnect_0:sgdma_rx_descriptor_read_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	wire  [31:0] sgdma_tx_descriptor_read_readdata;                          // mm_interconnect_0:sgdma_tx_descriptor_read_readdata -> sgdma_tx:descriptor_read_readdata
	wire         sgdma_tx_descriptor_read_waitrequest;                       // mm_interconnect_0:sgdma_tx_descriptor_read_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	wire  [31:0] sgdma_tx_descriptor_read_address;                           // sgdma_tx:descriptor_read_address -> mm_interconnect_0:sgdma_tx_descriptor_read_address
	wire         sgdma_tx_descriptor_read_read;                              // sgdma_tx:descriptor_read_read -> mm_interconnect_0:sgdma_tx_descriptor_read_read
	wire         sgdma_tx_descriptor_read_readdatavalid;                     // mm_interconnect_0:sgdma_tx_descriptor_read_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	wire         sgdma_rx_descriptor_write_waitrequest;                      // mm_interconnect_0:sgdma_rx_descriptor_write_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	wire  [31:0] sgdma_rx_descriptor_write_address;                          // sgdma_rx:descriptor_write_address -> mm_interconnect_0:sgdma_rx_descriptor_write_address
	wire         sgdma_rx_descriptor_write_write;                            // sgdma_rx:descriptor_write_write -> mm_interconnect_0:sgdma_rx_descriptor_write_write
	wire  [31:0] sgdma_rx_descriptor_write_writedata;                        // sgdma_rx:descriptor_write_writedata -> mm_interconnect_0:sgdma_rx_descriptor_write_writedata
	wire         sgdma_tx_descriptor_write_waitrequest;                      // mm_interconnect_0:sgdma_tx_descriptor_write_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	wire  [31:0] sgdma_tx_descriptor_write_address;                          // sgdma_tx:descriptor_write_address -> mm_interconnect_0:sgdma_tx_descriptor_write_address
	wire         sgdma_tx_descriptor_write_write;                            // sgdma_tx:descriptor_write_write -> mm_interconnect_0:sgdma_tx_descriptor_write_write
	wire  [31:0] sgdma_tx_descriptor_write_writedata;                        // sgdma_tx:descriptor_write_writedata -> mm_interconnect_0:sgdma_tx_descriptor_write_writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;     // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;  // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_tse_control_port_readdata;                // tse:reg_data_out -> mm_interconnect_0:tse_control_port_readdata
	wire         mm_interconnect_0_tse_control_port_waitrequest;             // tse:reg_busy -> mm_interconnect_0:tse_control_port_waitrequest
	wire   [7:0] mm_interconnect_0_tse_control_port_address;                 // mm_interconnect_0:tse_control_port_address -> tse:reg_addr
	wire         mm_interconnect_0_tse_control_port_read;                    // mm_interconnect_0:tse_control_port_read -> tse:reg_rd
	wire         mm_interconnect_0_tse_control_port_write;                   // mm_interconnect_0:tse_control_port_write -> tse:reg_wr
	wire  [31:0] mm_interconnect_0_tse_control_port_writedata;               // mm_interconnect_0:tse_control_port_writedata -> tse:reg_data_in
	wire         mm_interconnect_0_sgdma_rx_csr_chipselect;                  // mm_interconnect_0:sgdma_rx_csr_chipselect -> sgdma_rx:csr_chipselect
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_readdata;                    // sgdma_rx:csr_readdata -> mm_interconnect_0:sgdma_rx_csr_readdata
	wire   [3:0] mm_interconnect_0_sgdma_rx_csr_address;                     // mm_interconnect_0:sgdma_rx_csr_address -> sgdma_rx:csr_address
	wire         mm_interconnect_0_sgdma_rx_csr_read;                        // mm_interconnect_0:sgdma_rx_csr_read -> sgdma_rx:csr_read
	wire         mm_interconnect_0_sgdma_rx_csr_write;                       // mm_interconnect_0:sgdma_rx_csr_write -> sgdma_rx:csr_write
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_writedata;                   // mm_interconnect_0:sgdma_rx_csr_writedata -> sgdma_rx:csr_writedata
	wire         mm_interconnect_0_sgdma_tx_csr_chipselect;                  // mm_interconnect_0:sgdma_tx_csr_chipselect -> sgdma_tx:csr_chipselect
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_readdata;                    // sgdma_tx:csr_readdata -> mm_interconnect_0:sgdma_tx_csr_readdata
	wire   [3:0] mm_interconnect_0_sgdma_tx_csr_address;                     // mm_interconnect_0:sgdma_tx_csr_address -> sgdma_tx:csr_address
	wire         mm_interconnect_0_sgdma_tx_csr_read;                        // mm_interconnect_0:sgdma_tx_csr_read -> sgdma_tx:csr_read
	wire         mm_interconnect_0_sgdma_tx_csr_write;                       // mm_interconnect_0:sgdma_tx_csr_write -> sgdma_tx:csr_write
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_writedata;                   // mm_interconnect_0:sgdma_tx_csr_writedata -> sgdma_tx:csr_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;    // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest; // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_main_memory_s1_chipselect;                // mm_interconnect_0:main_memory_s1_chipselect -> main_memory:chipselect
	wire  [31:0] mm_interconnect_0_main_memory_s1_readdata;                  // main_memory:readdata -> mm_interconnect_0:main_memory_s1_readdata
	wire  [16:0] mm_interconnect_0_main_memory_s1_address;                   // mm_interconnect_0:main_memory_s1_address -> main_memory:address
	wire   [3:0] mm_interconnect_0_main_memory_s1_byteenable;                // mm_interconnect_0:main_memory_s1_byteenable -> main_memory:byteenable
	wire         mm_interconnect_0_main_memory_s1_write;                     // mm_interconnect_0:main_memory_s1_write -> main_memory:write
	wire  [31:0] mm_interconnect_0_main_memory_s1_writedata;                 // mm_interconnect_0:main_memory_s1_writedata -> main_memory:writedata
	wire         mm_interconnect_0_main_memory_s1_clken;                     // mm_interconnect_0:main_memory_s1_clken -> main_memory:clken
	wire         mm_interconnect_0_descriptor_memory_s1_chipselect;          // mm_interconnect_0:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_readdata;            // descriptor_memory:readdata -> mm_interconnect_0:descriptor_memory_s1_readdata
	wire   [9:0] mm_interconnect_0_descriptor_memory_s1_address;             // mm_interconnect_0:descriptor_memory_s1_address -> descriptor_memory:address
	wire   [3:0] mm_interconnect_0_descriptor_memory_s1_byteenable;          // mm_interconnect_0:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	wire         mm_interconnect_0_descriptor_memory_s1_write;               // mm_interconnect_0:descriptor_memory_s1_write -> descriptor_memory:write
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_writedata;           // mm_interconnect_0:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	wire         mm_interconnect_0_descriptor_memory_s1_clken;               // mm_interconnect_0:descriptor_memory_s1_clken -> descriptor_memory:clken
	wire         mm_interconnect_0_ram_block_s1_chipselect;                  // mm_interconnect_0:RAM_block_s1_chipselect -> RAM_block:chipselect
	wire  [31:0] mm_interconnect_0_ram_block_s1_readdata;                    // RAM_block:readdata -> mm_interconnect_0:RAM_block_s1_readdata
	wire   [9:0] mm_interconnect_0_ram_block_s1_address;                     // mm_interconnect_0:RAM_block_s1_address -> RAM_block:address
	wire   [3:0] mm_interconnect_0_ram_block_s1_byteenable;                  // mm_interconnect_0:RAM_block_s1_byteenable -> RAM_block:byteenable
	wire         mm_interconnect_0_ram_block_s1_write;                       // mm_interconnect_0:RAM_block_s1_write -> RAM_block:write
	wire  [31:0] mm_interconnect_0_ram_block_s1_writedata;                   // mm_interconnect_0:RAM_block_s1_writedata -> RAM_block:writedata
	wire         mm_interconnect_0_ram_block_s1_clken;                       // mm_interconnect_0:RAM_block_s1_clken -> RAM_block:clken
	wire         irq_mapper_receiver0_irq;                                   // sgdma_rx:csr_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                   // sgdma_tx:csr_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                   // ext_irq_adapter_0:interrupt_sender_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                   // jtag_uart:av_irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                       // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         tse_receive_valid;                                          // tse:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire  [31:0] tse_receive_data;                                           // tse:ff_rx_data -> avalon_st_adapter:in_0_data
	wire         tse_receive_ready;                                          // avalon_st_adapter:in_0_ready -> tse:ff_rx_rdy
	wire         tse_receive_startofpacket;                                  // tse:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire         tse_receive_endofpacket;                                    // tse:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire   [5:0] tse_receive_error;                                          // tse:rx_err -> avalon_st_adapter:in_0_error
	wire   [1:0] tse_receive_empty;                                          // tse:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                              // avalon_st_adapter:out_0_valid -> sgdma_rx:in_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                               // avalon_st_adapter:out_0_data -> sgdma_rx:in_data
	wire         avalon_st_adapter_out_0_ready;                              // sgdma_rx:in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                      // avalon_st_adapter:out_0_startofpacket -> sgdma_rx:in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                        // avalon_st_adapter:out_0_endofpacket -> sgdma_rx:in_endofpacket
	wire   [5:0] avalon_st_adapter_out_0_error;                              // avalon_st_adapter:out_0_error -> sgdma_rx:in_error
	wire   [1:0] avalon_st_adapter_out_0_empty;                              // avalon_st_adapter:out_0_empty -> sgdma_rx:in_empty
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [RAM_block:reset, avalon_st_adapter:in_rst_0_reset, descriptor_memory:reset, irq_mapper:reset, jtag_uart:rst_n, main_memory:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator:in_reset, sgdma_rx:system_reset_n, sgdma_tx:system_reset_n, tse:reset]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [RAM_block:reset_req, descriptor_memory:reset_req, main_memory:reset_req, nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                     // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> ext_irq_adapter_0:reset

	nios_system_RAM_block ram_block (
		.address     (mm_interconnect_0_ram_block_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_ram_block_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_ram_block_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_ram_block_s1_write),      //       .write
		.readdata    (mm_interconnect_0_ram_block_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_ram_block_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_ram_block_s1_byteenable), //       .byteenable
		.address2    (ram_block_s2_address),                      //     s2.address
		.chipselect2 (ram_block_s2_chipselect),                   //       .chipselect
		.clken2      (ram_block_s2_clken),                        //       .clken
		.write2      (ram_block_s2_write),                        //       .write
		.readdata2   (ram_block_s2_readdata),                     //       .readdata
		.writedata2  (ram_block_s2_writedata),                    //       .writedata
		.byteenable2 (ram_block_s2_byteenable),                   //       .byteenable
		.clk         (clk_clk),                                   //   clk1.clk
		.reset       (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),        //       .reset_req
		.freeze      (1'b0)                                       // (terminated)
	);

	nios_system_descriptor_memory descriptor_memory (
		.clk        (clk_clk),                                           //   clk1.clk
		.address    (mm_interconnect_0_descriptor_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_descriptor_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_descriptor_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_descriptor_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_descriptor_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_descriptor_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_descriptor_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                    // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),                //       .reset_req
		.freeze     (1'b0)                                               // (terminated)
	);

	ext_irq_adapter ext_irq_adapter_0 (
		.interrupt_sender_irq (irq_mapper_receiver2_irq),           // interrupt_sender.irq
		.irq_input            (ext_irq_adapter_new_signal),         //      conduit_end.new_signal
		.clk                  (clk_clk),                            //       clock_sink.clk
		.reset                (rst_controller_001_reset_out_reset)  //       reset_sink.reset
	);

	nios_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                   //               irq.irq
	);

	nios_system_main_memory main_memory (
		.clk        (clk_clk),                                     //   clk1.clk
		.address    (mm_interconnect_0_main_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_main_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_main_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_main_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_main_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_main_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_main_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze     (1'b0)                                         // (terminated)
	);

	nios_system_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	nios_system_sgdma_rx sgdma_rx (
		.clk                           (clk_clk),                                   //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),           //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_rx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_rx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_rx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_rx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_rx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_rx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_rx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_rx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_rx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_rx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),                  //          csr_irq.irq
		.in_startofpacket              (avalon_st_adapter_out_0_startofpacket),     //               in.startofpacket
		.in_endofpacket                (avalon_st_adapter_out_0_endofpacket),       //                 .endofpacket
		.in_data                       (avalon_st_adapter_out_0_data),              //                 .data
		.in_valid                      (avalon_st_adapter_out_0_valid),             //                 .valid
		.in_ready                      (avalon_st_adapter_out_0_ready),             //                 .ready
		.in_empty                      (avalon_st_adapter_out_0_empty),             //                 .empty
		.in_error                      (avalon_st_adapter_out_0_error),             //                 .error
		.m_write_waitrequest           (sgdma_rx_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (sgdma_rx_m_write_address),                  //                 .address
		.m_write_write                 (sgdma_rx_m_write_write),                    //                 .write
		.m_write_writedata             (sgdma_rx_m_write_writedata),                //                 .writedata
		.m_write_byteenable            (sgdma_rx_m_write_byteenable)                //                 .byteenable
	);

	nios_system_sgdma_tx sgdma_tx (
		.clk                           (clk_clk),                                   //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),           //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_tx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_tx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_tx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_tx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_tx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_tx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_tx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_tx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_tx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_tx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver1_irq),                  //          csr_irq.irq
		.m_read_readdata               (sgdma_tx_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_tx_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_tx_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_tx_m_read_read),                      //                 .read
		.out_data                      (sgdma_tx_out_data),                         //              out.data
		.out_valid                     (sgdma_tx_out_valid),                        //                 .valid
		.out_ready                     (sgdma_tx_out_ready),                        //                 .ready
		.out_endofpacket               (sgdma_tx_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (sgdma_tx_out_startofpacket),                //                 .startofpacket
		.out_empty                     (sgdma_tx_out_empty),                        //                 .empty
		.out_error                     (sgdma_tx_out_error)                         //                 .error
	);

	nios_system_tse tse (
		.clk           (clk_clk),                                        // control_port_clock_connection.clk
		.reset         (rst_controller_reset_out_reset),                 //              reset_connection.reset
		.reg_addr      (mm_interconnect_0_tse_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_0_tse_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_0_tse_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_0_tse_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_0_tse_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_0_tse_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (tse_pcs_mac_tx_clock_connection_clk),            //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (tse_pcs_mac_rx_clock_connection_clk),            //   pcs_mac_rx_clock_connection.clk
		.set_10        (tse_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (tse_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (tse_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (tse_mac_status_connection_ena_10),               //                              .ena_10
		.rgmii_in      (tse_mac_rgmii_connection_rgmii_in),              //          mac_rgmii_connection.rgmii_in
		.rgmii_out     (tse_mac_rgmii_connection_rgmii_out),             //                              .rgmii_out
		.rx_control    (tse_mac_rgmii_connection_rx_control),            //                              .rx_control
		.tx_control    (tse_mac_rgmii_connection_tx_control),            //                              .tx_control
		.ff_rx_clk     (clk_clk),                                        //      receive_clock_connection.clk
		.ff_tx_clk     (clk_clk),                                        //     transmit_clock_connection.clk
		.ff_rx_data    (tse_receive_data),                               //                       receive.data
		.ff_rx_eop     (tse_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (tse_receive_error),                              //                              .error
		.ff_rx_mod     (tse_receive_empty),                              //                              .empty
		.ff_rx_rdy     (tse_receive_ready),                              //                              .ready
		.ff_rx_sop     (tse_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (tse_receive_valid),                              //                              .valid
		.ff_tx_data    (sgdma_tx_out_data),                              //                      transmit.data
		.ff_tx_eop     (sgdma_tx_out_endofpacket),                       //                              .endofpacket
		.ff_tx_err     (sgdma_tx_out_error),                             //                              .error
		.ff_tx_mod     (sgdma_tx_out_empty),                             //                              .empty
		.ff_tx_rdy     (sgdma_tx_out_ready),                             //                              .ready
		.ff_tx_sop     (sgdma_tx_out_startofpacket),                     //                              .startofpacket
		.ff_tx_wren    (sgdma_tx_out_valid),                             //                              .valid
		.mdc           (tse_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in       (tse_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out      (tse_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen      (tse_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.magic_wakeup  (),                                               //           mac_misc_connection.magic_wakeup
		.magic_sleep_n (),                                               //                              .magic_sleep_n
		.ff_tx_crc_fwd (),                                               //                              .ff_tx_crc_fwd
		.ff_tx_septy   (),                                               //                              .ff_tx_septy
		.tx_ff_uflow   (),                                               //                              .tx_ff_uflow
		.ff_tx_a_full  (),                                               //                              .ff_tx_a_full
		.ff_tx_a_empty (),                                               //                              .ff_tx_a_empty
		.rx_err_stat   (),                                               //                              .rx_err_stat
		.rx_frm_type   (),                                               //                              .rx_frm_type
		.ff_rx_dsav    (),                                               //                              .ff_rx_dsav
		.ff_rx_a_full  (),                                               //                              .ff_rx_a_full
		.ff_rx_a_empty ()                                                //                              .ff_rx_a_empty
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.sys_clk_clk_clk                                (clk_clk),                                                    //                              sys_clk_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                           //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                       //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                        //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                              //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                          //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                             //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                         //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                       //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                    //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                       //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                   //                                         .readdata
		.sgdma_rx_descriptor_read_address               (sgdma_rx_descriptor_read_address),                           //                 sgdma_rx_descriptor_read.address
		.sgdma_rx_descriptor_read_waitrequest           (sgdma_rx_descriptor_read_waitrequest),                       //                                         .waitrequest
		.sgdma_rx_descriptor_read_read                  (sgdma_rx_descriptor_read_read),                              //                                         .read
		.sgdma_rx_descriptor_read_readdata              (sgdma_rx_descriptor_read_readdata),                          //                                         .readdata
		.sgdma_rx_descriptor_read_readdatavalid         (sgdma_rx_descriptor_read_readdatavalid),                     //                                         .readdatavalid
		.sgdma_rx_descriptor_write_address              (sgdma_rx_descriptor_write_address),                          //                sgdma_rx_descriptor_write.address
		.sgdma_rx_descriptor_write_waitrequest          (sgdma_rx_descriptor_write_waitrequest),                      //                                         .waitrequest
		.sgdma_rx_descriptor_write_write                (sgdma_rx_descriptor_write_write),                            //                                         .write
		.sgdma_rx_descriptor_write_writedata            (sgdma_rx_descriptor_write_writedata),                        //                                         .writedata
		.sgdma_rx_m_write_address                       (sgdma_rx_m_write_address),                                   //                         sgdma_rx_m_write.address
		.sgdma_rx_m_write_waitrequest                   (sgdma_rx_m_write_waitrequest),                               //                                         .waitrequest
		.sgdma_rx_m_write_byteenable                    (sgdma_rx_m_write_byteenable),                                //                                         .byteenable
		.sgdma_rx_m_write_write                         (sgdma_rx_m_write_write),                                     //                                         .write
		.sgdma_rx_m_write_writedata                     (sgdma_rx_m_write_writedata),                                 //                                         .writedata
		.sgdma_tx_descriptor_read_address               (sgdma_tx_descriptor_read_address),                           //                 sgdma_tx_descriptor_read.address
		.sgdma_tx_descriptor_read_waitrequest           (sgdma_tx_descriptor_read_waitrequest),                       //                                         .waitrequest
		.sgdma_tx_descriptor_read_read                  (sgdma_tx_descriptor_read_read),                              //                                         .read
		.sgdma_tx_descriptor_read_readdata              (sgdma_tx_descriptor_read_readdata),                          //                                         .readdata
		.sgdma_tx_descriptor_read_readdatavalid         (sgdma_tx_descriptor_read_readdatavalid),                     //                                         .readdatavalid
		.sgdma_tx_descriptor_write_address              (sgdma_tx_descriptor_write_address),                          //                sgdma_tx_descriptor_write.address
		.sgdma_tx_descriptor_write_waitrequest          (sgdma_tx_descriptor_write_waitrequest),                      //                                         .waitrequest
		.sgdma_tx_descriptor_write_write                (sgdma_tx_descriptor_write_write),                            //                                         .write
		.sgdma_tx_descriptor_write_writedata            (sgdma_tx_descriptor_write_writedata),                        //                                         .writedata
		.sgdma_tx_m_read_address                        (sgdma_tx_m_read_address),                                    //                          sgdma_tx_m_read.address
		.sgdma_tx_m_read_waitrequest                    (sgdma_tx_m_read_waitrequest),                                //                                         .waitrequest
		.sgdma_tx_m_read_read                           (sgdma_tx_m_read_read),                                       //                                         .read
		.sgdma_tx_m_read_readdata                       (sgdma_tx_m_read_readdata),                                   //                                         .readdata
		.sgdma_tx_m_read_readdatavalid                  (sgdma_tx_m_read_readdatavalid),                              //                                         .readdatavalid
		.descriptor_memory_s1_address                   (mm_interconnect_0_descriptor_memory_s1_address),             //                     descriptor_memory_s1.address
		.descriptor_memory_s1_write                     (mm_interconnect_0_descriptor_memory_s1_write),               //                                         .write
		.descriptor_memory_s1_readdata                  (mm_interconnect_0_descriptor_memory_s1_readdata),            //                                         .readdata
		.descriptor_memory_s1_writedata                 (mm_interconnect_0_descriptor_memory_s1_writedata),           //                                         .writedata
		.descriptor_memory_s1_byteenable                (mm_interconnect_0_descriptor_memory_s1_byteenable),          //                                         .byteenable
		.descriptor_memory_s1_chipselect                (mm_interconnect_0_descriptor_memory_s1_chipselect),          //                                         .chipselect
		.descriptor_memory_s1_clken                     (mm_interconnect_0_descriptor_memory_s1_clken),               //                                         .clken
		.jtag_uart_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),      //              jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),        //                                         .write
		.jtag_uart_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),         //                                         .read
		.jtag_uart_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),     //                                         .readdata
		.jtag_uart_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),    //                                         .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),  //                                         .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),   //                                         .chipselect
		.main_memory_s1_address                         (mm_interconnect_0_main_memory_s1_address),                   //                           main_memory_s1.address
		.main_memory_s1_write                           (mm_interconnect_0_main_memory_s1_write),                     //                                         .write
		.main_memory_s1_readdata                        (mm_interconnect_0_main_memory_s1_readdata),                  //                                         .readdata
		.main_memory_s1_writedata                       (mm_interconnect_0_main_memory_s1_writedata),                 //                                         .writedata
		.main_memory_s1_byteenable                      (mm_interconnect_0_main_memory_s1_byteenable),                //                                         .byteenable
		.main_memory_s1_chipselect                      (mm_interconnect_0_main_memory_s1_chipselect),                //                                         .chipselect
		.main_memory_s1_clken                           (mm_interconnect_0_main_memory_s1_clken),                     //                                         .clken
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                         .debugaccess
		.RAM_block_s1_address                           (mm_interconnect_0_ram_block_s1_address),                     //                             RAM_block_s1.address
		.RAM_block_s1_write                             (mm_interconnect_0_ram_block_s1_write),                       //                                         .write
		.RAM_block_s1_readdata                          (mm_interconnect_0_ram_block_s1_readdata),                    //                                         .readdata
		.RAM_block_s1_writedata                         (mm_interconnect_0_ram_block_s1_writedata),                   //                                         .writedata
		.RAM_block_s1_byteenable                        (mm_interconnect_0_ram_block_s1_byteenable),                  //                                         .byteenable
		.RAM_block_s1_chipselect                        (mm_interconnect_0_ram_block_s1_chipselect),                  //                                         .chipselect
		.RAM_block_s1_clken                             (mm_interconnect_0_ram_block_s1_clken),                       //                                         .clken
		.sgdma_rx_csr_address                           (mm_interconnect_0_sgdma_rx_csr_address),                     //                             sgdma_rx_csr.address
		.sgdma_rx_csr_write                             (mm_interconnect_0_sgdma_rx_csr_write),                       //                                         .write
		.sgdma_rx_csr_read                              (mm_interconnect_0_sgdma_rx_csr_read),                        //                                         .read
		.sgdma_rx_csr_readdata                          (mm_interconnect_0_sgdma_rx_csr_readdata),                    //                                         .readdata
		.sgdma_rx_csr_writedata                         (mm_interconnect_0_sgdma_rx_csr_writedata),                   //                                         .writedata
		.sgdma_rx_csr_chipselect                        (mm_interconnect_0_sgdma_rx_csr_chipselect),                  //                                         .chipselect
		.sgdma_tx_csr_address                           (mm_interconnect_0_sgdma_tx_csr_address),                     //                             sgdma_tx_csr.address
		.sgdma_tx_csr_write                             (mm_interconnect_0_sgdma_tx_csr_write),                       //                                         .write
		.sgdma_tx_csr_read                              (mm_interconnect_0_sgdma_tx_csr_read),                        //                                         .read
		.sgdma_tx_csr_readdata                          (mm_interconnect_0_sgdma_tx_csr_readdata),                    //                                         .readdata
		.sgdma_tx_csr_writedata                         (mm_interconnect_0_sgdma_tx_csr_writedata),                   //                                         .writedata
		.sgdma_tx_csr_chipselect                        (mm_interconnect_0_sgdma_tx_csr_chipselect),                  //                                         .chipselect
		.tse_control_port_address                       (mm_interconnect_0_tse_control_port_address),                 //                         tse_control_port.address
		.tse_control_port_write                         (mm_interconnect_0_tse_control_port_write),                   //                                         .write
		.tse_control_port_read                          (mm_interconnect_0_tse_control_port_read),                    //                                         .read
		.tse_control_port_readdata                      (mm_interconnect_0_tse_control_port_readdata),                //                                         .readdata
		.tse_control_port_writedata                     (mm_interconnect_0_tse_control_port_writedata),               //                                         .writedata
		.tse_control_port_waitrequest                   (mm_interconnect_0_tse_control_port_waitrequest)              //                                         .waitrequest
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	nios_system_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (6),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                               // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (tse_receive_data),                      //     in_0.data
		.in_0_valid          (tse_receive_valid),                     //         .valid
		.in_0_ready          (tse_receive_ready),                     //         .ready
		.in_0_startofpacket  (tse_receive_startofpacket),             //         .startofpacket
		.in_0_endofpacket    (tse_receive_endofpacket),               //         .endofpacket
		.in_0_empty          (tse_receive_empty),                     //         .empty
		.in_0_error          (tse_receive_error),                     //         .error
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (),                                       //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
