��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?������e�eZԒ��;����d�gbKK��V�ƪ9w)�32��:eig(�)divIc�I�����"�9��,���I1�
p��?ᑽ��a�of�ҥ@
��f������=��䪿�8����1�K�J٥ǆ�����mHkS�h��]�����=Ï�L�%�-&SUf|gt�t�#�Գ
�c��AP���������D�8��{���	+q�9 ��T��B�3=�H�|E��td���"�&�����V��2�|���	�ݙQ��Q�fpf2����Y�����Kt�>!�ߔ�`��7��&}u ���|l��k�����l�����'R�1�+�4��V�֮@���%��yy��U�qA8#%�y�c��_�ޔuШ率���I���t�w��b����:����
��ǄJ�qf��G@r6@�$�:�V��Px�C}ݼ�A*�(X���`�7�:A��kN�$M���������k���E9�2J{۠~�؏�ms�RH��Er��5j�G�3���w���m�xt�Te}vMu��7B�������0,�����_r�ꈳgy��':�A�LyS �̱���9�c���Dޚ��Mc����=�>��F:�� �"r���f_�R��k>]B$�~2��ݕx�f���8B�&^BLe�y��<�z���#ЯS_o.��Z�ר��eQ�#?'�ݼ�t�$�y�n��+}��A Li�X`�r�u����6���B���̘h')�#�K��VB[��/�.?fv [Lz����6��g>?ő;N~������wt��>4�A�f���!>��W�	��k|��Z��\�3WA���/O�Y�a�A[�ݞ�G��+?!9 .�!��!�'P.G� )5%�B�$HxijFo$�L�N�η���Ŵ�0Xd�|�tE�|&[O�~��Q}=�2�x!��XW��N*I�+���������<O���n|�1X%�3�K��X�x�y\�v��BJ�����'o�q�6�6_E:F~)!���J��y�
�~�V�k��%{�v�M����]��V+�7v1Σ���֧s�Q��L^;�̌d�����u���ǏxYm��v(`*���rj�"
�sa�((\ZTі��b�/�f//o��6G��\pl��J�Q�'�$�tM�V�S�7�"�h���64�!���KE!������Ỳ�G%z�>s�%�%�-x�Q*ӒB\�<�+����V����O.^�bӓ��sƱ��3����������*NһM�W�)�5r���=�zH�JN_��,�e��b�ʨ�<��=/�%��+�3 ����;j&
q���X���K8@�Hz��t����r��J����ڝ)}D)Õ7��(#��M$Ԅ��B�����h��Xq�KЮZ"����E�/%�N/�U�Y����>E�jy�+*�X8��.t��r �ч�Y��"��a,���ĵN���N���^;]�4���j@�k�s��M
�Z?W.GB��zK�)��t���#������,(��Y�&��sY�>��'�)�'B�]�@�z��%�O�C�Ser��g��44pG��<V�`�{���(ْ7L��#�S3�($�V����pq���Y3 ��c��l|�HaG��->�n �k��yX���7����)0���e�ɯ�<��׫�
���P~�q9Bq��]���\���=l<y�]�*��HQ���bX��c��|�b���o�Fs"a 1J�q*�s«�Q�B޵ukn��pr�MPE�)�l���f�c��k~�_Y770�x�  p�֞�*�D���A�H5��o�0��f����g2S�.��+Ce��p�&�{���0悖S�eDMɻ,�К6<�>��3^E\��þ*B���hC��I��8�5��`�k�ǐ@g ~̭�W�d/$�A��r1k�6B�1x8�y���c@.okv-�!�y`���|�;_9�x��b�?����x�j����m֒���λ޺�#�&��4X�dπ�f�xI�M����!-=:-�M��d@����D��8�%9ҟ�����V��	�n涑J��)�����s�r��N�e�mkT����)U����Qf�p$�JS�Y�ߦ2`��|��v�5BT�l~_{�q�t�h��N�vz�|rE����P�'�i�
)�YՐ�yɼcfq��!��R$ۼy劍��V\��ϴ7�+��ءA�+��fc��d��+u�/�1u(�)�m��d&�?��ЃT��wq���i-OޠW6��e�iNV��R�]<�L��Akh$����^�I�[�> �۠�"z.�,�N��.<k�P^p)Y��}d���˳E1-R!i��w���,��n�i�����MI���giG�^�t�"7�4�_�_��q��쒴o`摣YJ��6Q��S��7�'��� v�b�3qҡ��^JR���Ǎ�¤�E%oLY�ګC�x$0�&p�RBEuF�YڭL�&��E+���[��Y©�����q �^�%��\�����Q�Dۡ�qN�I#�9��	�C�z����*�9���i���!=eͲ4$/��p�O����E+�R��}_�}��D��'
Ϝ���&�ZQe���+��Z<���'����� �`>W�ˊnxa$c���d��om8.���N�=
'і\�3���l�ӫN�������6���KKn�?^ߪ1��J|s)��$9��LQ;���V&��'}G*�����D�_�~�`w��R�����'ȟ��憽�~,M�YvJl$j _�b����r�$��,_g�g&餿��*0bV-_� j�o Ϳ&μ
�ۀ��X���ݵ�q*&�kL"Zs�z-
����/S����$�:me�4��˚N��^���:����u��6��~qܼ �j!���C�3Dϸ�9���]�e���ۃ�f����6��53���
Z�a�PU}�4I�?�+���X�ރ�F����SP�v�Y;�zw{x�����'��>n���k�3���$�O���x��6���a�c9(O�AQL��`9�+���$S�y�9L�QĲ���9��X�EȢ����B��]�Ǩ �c�
�L��2�UL�@�y�*��1�^�y�{���/�k�X��Z������a�ݰ%~�֠�`�b	l]�)jz`�j�nAg���\��5��2��b�M��B�࿰;Na��O��n�AS�b�����N���Fo�N�6z4�{�xů�D��G\�pc��l��1"���)TƓ�\�^�*܊��O�d9�=i�t�A �E�V���nM<��H�;��d`)HS�Z�R����x�^��y���ʿ�H���;Y�����u��!Y��Q��{������0�wĤ�Ғ?�5W�u	B6H�Xd��S�':a���ß����>���W�s	����c,-�L�<��&�������=�y����_�mRA�P�[��-��});�
ة��ٱ��=|�r�����Iy{��㳉�� ɛ����� �,�u�?	�U����6��)g���_�ʡ����B@,}f�o�a?�?�Y�E�&�io���$WA��(!�]��t�:�ٻ�!����EK�}O�͊�A�����i!�7���"K�]A���a�tO=�W���9�W���lu}pkȼ���Sl����'^&G~�׭��3�谻�X�;yŖ|�;-'<�Z�j���}�*@w�	�+
�:(�,a9��[��&�����A�oN��j����l�X0[��:BJB�:���G�Kڽx���L$���lk���G���� SU���Ix(\v�:���G��m�%o[�^o�>�S9Tn��(�?��ןh����!�^z{�����@ٳ�y�����eƶ�������b5N
�j��E�Դ����!�`�����A�)WH��p ������0n�ZsR�� �1�ڊ�uhM�V:�z.a�.:֠��ܰ4 �Y�/$��e��1q�P��6`���[�C63����d �9��>!��0�mc1t�a{��:��pO���>��>h�M��k&��m��-�b<h��^��Ӹ�T������<��uM�3�M��H�I���U0�ߝ��=�{Μ��6��M]��?e���yR�G+��M����G$mHyU,<8�~ys�ۋ�[��Gr��Ɣ�nb��a}�Z�H㟆b�����$~ZO����g@��\G@�K�j�w����b�S�낕�m���呑_x���߭��e��WH���\�
�i�{��%ȣ��@�ʽ�Z�J;24���%W�P)c_���c�H�td�|�3�