��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��yX(�C¥Jd(LR��h�Q�Xd�H��b'��� j�G2��Y�`/�YR-�r��Q�M���l-ý�b2 �P2�;�k�(M���*y��r=$���D��o8p�_i׊�ۓ2���⯚y9r�2A�I����O��9��p��\t��
uV߫���͠�:���%� ���3'����FK�uf�Z��f��  u|��̱�/	C��Il4B;�ycu2�I��ٌzǼ�U�m9��,�q���'0eת_!��QFhc:�"*�cIQ�$�^�E�dV�Bz���S��ǟW�@44�#��[�j)�:GI�i�܉n�&7���+�:;	Ӫ���1�d�	Y���G�$�Ҩk��s���Lw։:�B*�Rl���I|�eN��6;���:�ή%��B��n��ͳOL���̱�u8B��=�&�Uz�r�M��Y���M;��9�k����	e�h�:��[b�=	B(��󲂇�����i�ڞa�܅.G�����m4b/����	��q���9V\�I��E㫨�258�8T����ҝ�)�{Z�u3
k^�F'�rRE{Q�����I�X7w��"�rޠO
����L��|)��t���.��CŦ��/\r?��n�|����[�;����nY��	�k��\l��j��+�)�tX�'���;��|�<4��v�3�ƑF�!q�r����v�+L�� )�D#�1?���S�u���wu��m�IU�?��h�ۿcrM���+��un]�������l�Zg�/]6Wi$�)��U��۱��i�<_J��ߍw�I���G�0�߫���������x����쿇V"	�Q3�*_ �wc�<�����;�˵�[�E�m�Ba�J7��ʢ����������`�cЕ��]>���Yh��Kj��~��h��$�Q?��7dZ�;�bl_�u1u]�T�]�m��ų]��4���vMȱy 6ҳe=t��[}ɯ�,�,��)#IJ�=��<L�Hs�����ٓ�v���6 �]�� �<��~qR��H�*F˓x���VSS�gR�2K��O��H�50t���51ET#[��)ٖ���8���L@G����L$2�E4��2�s.F03m�;�[�ԏY1�G�[���f3k_�Ll��R/5�i�'g]&��g�g�<j+z�E�W� �(�D���װ�<�@��@O���	��H���4���R1�R�*;�h>���j�|~�;v�q%���"��Ѭ <���62���?4���G�|�rCYЦ�4�y��o3�'+�<}���j��nS��L#�(��9�=�_�2�kn��Px2;�BBQ��q�i=�F�J]Is��z+�bh�1�C_
��=����o�&�,bͅ�z��'<��@�O=�	"h��E�e� ��TYh�Í4lX������_�,)����%x��z�zPV���5��^��D@�ܗK>���Q9:�C���x�+��T���uR':�Y��h�����w���X�fi��1��Sʣ��E�+��ݐ��L��4���v�,/�:.�C�O�;VT��Z�9��ؗ�421���EbfM��O���'o䂼/�<׉��c�(�^\�4��˛w�:.j�K��0*�?r޼��&m�c8 �y���Ԍ�a����5�\>c}�i@4Ar�H	
��g�_�܈i@���z����z�syz���88U��٫�3��1UT���9�R�V���G(��H]T{[��>�����T�A0eZRq��V�F���Q��;����ڒҗ0����ϗ� ǣ�3���Z���Զ0&:w����dc�E�.TO)���K�
�`����5us��,�K5�*����0��տ���}�)��f�L�K� T��J�a'365��$s ӽ���A���
�b����d~�BD/9��DR��m�%�p@��X���Ȝ�d��6�f*7h�X�4Bg;NY=�/�����P4ʃ����B?SDU�|t�FG(A˫=�����R�����9e�t�0%��]�٠u[~���?"��~'"<�-�̠$'�3K�y��`�t�^iT���\%y*F��k�����&�o)��b��Ix�<*�+܅��)N��a��_�
��L��%�4ł��q�Є���$�Tm�6d1=��5�j�AOm�4���ػ;#7�k���'k��+
k��2�� �=�9��s�#�|�Ip�(�t�-l����n �6a�o�|��ibҢ�La6����U�����%�� v���A�u#6Ů߫#b�m9�4�:/�C~��!��*���J��HC����⏀������yO�����py��_��A:��FH�R����{����+��"F��Ay�X���+�لP��7��-J�T�[1t��{� ��H�xظn��nC\�h���W|���H0h�S���kd����@w$���)��׌5d��4�E���0�o}#��V�d�����	b��܏ Y	wV�]��XvL�W/� �+��J�LL4i#t��,i���{�Ǭ�SEď��g[-@���c��@[�K3�t����+�G���i^ݩO	��_Î�/;��F�d�>����8�r�_�f���!�Ɑj�R4_�L*�q�A66�WFh\�bz��8��:�����Y�,O��d˖���}Qx �}@�N�#��h��6�WC �Gy1�}Nv�2�S<7t�>�><+o�P���^�%J�A@[�I�	.Sڐ���b����b���P孒K��WV
ml_%~�R��$x��F 8}��?1�jS�W8Ny;s�6�: ܚ�رI: �3��jYSKƮw�FM��O�B���J��⨿A�I�[d�
�HĊ���2����\]�rnV�,����t�I�Xߴ�+�����{.�"D��!!r!�UdL�^&��^ ds���ɲ��@E�AE�	�p�'a�O��}���#�|��7!~�wF<�OQ�6��NpMYd�]�^�è����Z�F�WAcF�w!Y3Ví�2�nH1��oypi'А�0����aw��2�w$V��"WW�?���W8�h,�g�5�ǃ*�aeN���^5AZ\m�c��T<nfY�|����\F�I����L�������7L|C$�*��Ӕ)i/`J ���"ne�����񁵦���g�K� �A ��z~�{�9��l�.^8�N�&T�4���X�?1�t)}wG�!!OИ5��W����"۪����t���U)�9!쨡>ϳ�e�~`/�>��$�# �G9�;�����~�H��m���T̮�ϣ���v�8�	ߟx����qX2"S�oܭ�gLۮ�o���H�p(�?8$����Y��'�H�r�D�����\���ni�I��ija�+
��O�)�Ԧ�P������u�a�L}YT���#$`\J�UͥՀ�UoL����H�N%	&���q҃�_�29�z)�a��`�7=��$ri��0$��jA�)O�p�������Z����*��9�����[0H����q��NY��ݪ4�CK�N�E��O�6�N�]�E�����=2ϛ��0��$VN�j1���N+�@�	�}O�|�g0� ��dZ���!�n�$0J(CnfR		��|�%�G8_)�6H	
��9�Clx9X)9}�q����0ɕ�o����G����Gu�"j��Y\�V�Y/�����`�П��+ �3�E��i�(�,�t�@l�sa�,��]�>I�F���FZ�3�*]UE�,]c����r!�@Z�UQ$�*�Uf��we"�Ԛ�*�y�4`��)�h�X��n����T`y�!b����Хn��o�%��wӮ�����Qhc�й����|�b���w�K�bI����j�O�!������	\�A�OM-z�TuZ�,3��-4hE_�{L���m�h��C�u�Ao��KK��tz`����mw�0���4\j ؙ�m#1�aqb�㨻��s;��=Tj�r�!+5�[�\�=�Z�⿹�Z_��}��3�����ʇ�'R��w�cc�"� ��A��?J=�xc�qB40��t-�l^kz<x�:!�@����:����h�Ed$Q\G<8N� �%����7���T���n�:1��&�QADq�X<?�#�>1�9�=ƐJ�����DəWr$�h%o��_FY�cB�������u���8��j�a���.G�X{�� �l��ء��H���󙊪5Ϟ7t�nE{2�L�Gb]a��9��u*�+1O<c�s��s��S�	�Y^W&��7(�Wu��BD��¯4SO�
j["4U�D�]��lnm(���q?�<���x ؃b#��t����yLFd����x��5)�q�+���(�@�Q��8 u�����W�֣G�4�1�d?ڃUAC|ǃG3Da� �Q$�C�
��	�Fo�qY�p�9C�\o$#Sj�ih�K{��Ajm���R"[vu�o9I�i0KZ5r��Zv�B��3��DS��S/a}I@�Ҙ��[��R�		��7�!zS���0�e��$����g�M	B���MI����n9�:�P�6�!��V�1�YY��.?1�W���\���-{��)ψ�xE͞�S84�|��dH�� ��	�]�;����v��Cq]� �i�I���t+��.樎�*%v�'N�ǘ� dC<΍�T�bMm�1N���ui%�^-��?�>P�d�I ��ͱb쐍v�.^�=r@b̟�f���S��̇�$x6��0�@��v���x��_Hy�豭��=m�^��}�%b�T	͑����;A�'2�K" �Vysh����B�ꅜ}�5��zpL�#t��rVe���*�� ��j�i���t�쾍���ģ�b�Y�د�;Z;^~�Qc�lZ�ɳ�ݛ�}�n�t$>��T�6��$;�w?�о�xo�J�Y�����u�����ߦߍG;��x"����L�h��T=R�����(]�"-܂���j�M\�d�k����x�,|С���K/����{��ڣ]�8X>Үr�I������ ��9�b#��Rt�ͷ��$��y�����w�R��"��n����A	'�����Ri��2�������u[,��[���3���! yb��
�u	v�u�!3�[9�s��9B����_��Q$k3t;�z�����C壔o7(���T��W�L_����J�
d�J�5��Sc�a�6�h�X����QȈ�t��A��<�;�v^cn����DZ��j���zV�ii� I��yUAJy�@��{�Ž���l.�<Ӏ�[K	Wl�#��Kǟ�(�i�F��B`و��$v���ҍ_6N2�h�uJ�9�tWZJ~�c<y�D�����^x�}�rI3�]���!�ƺX��#�GW,�Vm,�j����[��*�L�d$�*U���U[1{M���'�*i�Ѡ:�ɹU>�Y?������CL��p_�!�T*g�>]��N��0'H�W�;X=د�y	<�(�5�D�%+���r�s�>�d9w~�-�r;Nvl��1�9g���W�F��%O�����ÏC�0��H�ۉ���7+��猇�G���H:��L����X�-�-�5�W��k@LY5�	>��[l-�~x�B��UmH`uC�U��=}bD�C�]���4�⊋짠Ӣ�i���K,Ю��:��[SA�)@��f�ڕ�d��k_���m[d;��F�,S�sa�v4�V54.#Rx,�/B���<JȮ��$!��BtA�����Nr��G��C`�}�-3�z���M��pB���tq;(�~���ά���j�\c|�t⯮��ة�S�4���1�M��.\(T�!�������s/K��ó��X����mz���o�U�!����cE��H�%ʥ��-�S��Z"%oo͍�͸a������'uiT�l&�/3?���,�$B�O�?����))b��޴���1\�w�C�3�uct�SbGdTaOĜ+b~hᮻ��u}R?2��I=���sL�%@�p���(Z(F��R��ɖ�����YYˏ�&l4���職#��Mbg=+AU����,	J���7!}��M�g.�get���B���?�^��������̛+�S�V~�V��ZQ�b��<��@N�(0t6�(�_gE�tT:�E� ��	'=9���;������� J��5}J��y�4;��ӱ1$�����Ѐ^73�������Z1�^2̽#F�7��s�7�Y�� ��i���X[X#?{��Vt�ˢ"Y%�GՌ>|��<eY?����_�y���&0,��*"-��R8��1f�>�P���;�!���@oX�s�\��q��=c?��><9h�{�=� W�VZ����ۗH̟�v���幇��jF⭮T������3�2=�� ��17�K%�t>rEU�;�k|l(��,���9v�-�W�%
W*�v�xY1���[f��y���Y�E��S�7�Ymb�>WJ�-	a��x~3A���Q�?��-ت�wJ�Ch`�n���j����g~Xrv[���7���D|H���|��+K#��[@�<Å�V<���3Aq���(s�>ɻ�R�q�C�)f�}�0�E�Xz������K:A�6 �1T��ӆ��\�lDIF�39[{�i���(�J9��?�����t�r�o%���Jڒ�N�!��h0F���