// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:14 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b5jljYzOCZfnQeO27vDwz8GQeSEh+I9CRIj6e/uoKC1T2gyUlVi5XzdkFFSrICfD
uZHdEjeC2X5nr1Fafgi+d5tF1QRBWe7G+0JD6mRtugbf0JzvK4NUfaXgLHlWTE4t
gOvv7InO7hk7xUU5tOKsXUK7cdsmvR70UkFedFVANnA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22912)
o/yQXdvwnfExuI8DY21weVwseWYkvUTkiH/fLo7ZHKh44+Auwtku1zhonFgQRaI8
Gmn4Yqxd+t+m0+1SEnmsUFkJSsv5OYAmIyj6bkxzoHHKgw5pxOJO/JFLUv/Pl1bE
nh9ErbSvHV7nJEYKuSYXg+fEzuIXdRX3DC0eI38onqOtn4oIxTU6WH5+YCf89fic
8cHYLsPFssoaciNFqYUuqxqNqjEVgdz9csOZRtNPM4btF+VzfuDGANTMiD759FZt
mUhnoraEH+N4CiRgfYXvsrx/Tzl8uPLwnWJl8sV+ieumRHu0Afr+9XU3qTJyU8/K
TPrz7+KQRJAPgMhxR2g7TN3+PzCjGQ5pws9qXFxfkmkbr5ApB2OBnmHeLrtVgDHa
MYLXK2pZVXo4XKurDXz+Wq9Q7HC5WRGjl+Kj+GJPPvkhtaYviQ4bF9B4jpXej+fb
xDLmuEfop/33UfxnMdlS/AfZp4p3eMp1moxdFlGuYcr8LnnI2WjURxTFZ4J7tOaI
GZhnXUugHo135N4ysYsPZtj/cwJ0Pv3EGFiHUcFi244Rv+qokcxIJzjhUmTyUXCh
zBhtYG7MFLlJ0/8sIXTkUxV5FI/qaL46tdUD0esN98ltbohNFrW4EjAMQd5S69Dz
gvEgwazE4oBJEaUL/xUBTy/jNJIxICy1avR0NMXT1P+B3NOWQhqSQS8NDXsAgqgz
eLsw0Rm/PuJcZnpnuT9Wbc5mmMz24a2Jc2Utusda9KM9suieY3Q5zjfcSx7TjHbg
+WPB4a55qmH9ftw9qSnby7/2NbABY/43X2x6Gddfi41Aq1fPGNho0g+uP7DYei2w
L+OqmE7c1nWQAqE1dLevrJQrsEWJKL83GlwrEsZfXTf6cFZ3XUbaAONPEhVYdRtc
3hDlH3s4aU85SIz8o57Qm/BCX5C8rQuhR/GaV5TY9h9s9lgQYtjxSrpxm7KbBl8h
h2EZPpCcbEnG4w8D//3bp+1vEjHAhZEOCbcn+MiA9yFST8nRVZ83KYF0gyESe9zG
I+DSTSdHRTNnPFPyOhWBWnUD/MEbeRL4P1a+//xDpGqdboDeFNnZAUMWxTXG6gyl
hNk+e1t/Y6TDNDrE8KLH/L/+Ia6O7MVaUIBwTPbOQ7ANaQKHDT1iH5Adc5nCGHaO
mLodmFEzL//HUDfYJH4b6pANpkaPJSR44vX0q7SX82Ca3ww25YliwZ4/CYJzzU/n
YnLseqZ7uNVnqFESEsXxzOqhjysMa/RpsyqFCZX3/FhPSZOEQkwecdAVQikU40OK
UlTqNE4C0eOwyUPU5g7aDeWmGbdTsLQYRqCpcZiZa/1NpkMhswmnUOTJGur2YZTw
vPCM8Dgq+u54/BlJ3doNYZVJr5vwdq8G87ZHWeF0Mp1p8WPGDNQhXG+f+GyAeqla
XVUtNHroc/uISBdzjhkc9TH4N7/zHdTJrh3Dcd6j9ngwgX6VFi98NTz1LvAQF4JM
AENFb0hiOrcEpAUgcZOu50Rpnar9m8eyahTmGGn8UtcBZXxDcSwljZOrwC8ziDdP
XPbHxQ9VWL8F8DGeEuXdWKsb+WozMdjpjrNuxNDyIJU/UXzMY6ZNlsFu+5wwdjI4
p6NC0FNpU9lyLxmAakBfeO1HyZqpYV63Aag0NSPlNWAEraSrutfjL0j6oKTYMddH
tb3giQGKZOO9AttkD/DXhVBNESMfzj56ZOG9PzOyj6UriiK+8jmtfe4jme8iE//W
FuaezNwu9gwUoEtFrJXEgkI5L+wgemoXuyyAgfqcQuv9yRgBXLqJFYEESor/KV1g
t8mYF27UAjx+cjmL06Yq+qz6rancxgmxLZo+wb03Opkgvkgx/ztHASWG06/iGq7f
WJ0xXoith1pF7yF25YxkGRbMt3b+8sb0ecWY6xLXrnRoTHqSlv50ewyroepQAPye
nrv9ntP63XeReGqdBIskAKzIGJxAyEX6FCFDkN7nM9n5Dy8F1fYaSkLkv/QpV+NF
iMojJk9BGufrEewqth5HKcxDyVMhFwtLBreAnfkHTmsIbF+kD13T72/QAwpYe+06
JlXgauFFgMabeyzBziSFB1SNjEVxBrfDYulbHrxDVUd6YJuHRUCcZoEhKhVauBbt
eB1aXdwq6d/MxmK9mDVx+X0qeY43k/pqr5NnXn522worSId+BLsgF5biIhc9llmJ
DcM1AinBAaCl4eqc0b47DqLjLdKgvCVLH0NcDfRqAERzxx2nNuEJJW4Xz3cVlJa8
q0qYx8qTqLhATmKG2fi6N/8SGgH4jzwWYfR85MPJz1n33dcjUR8G5ZBS0QTIFgbO
SkbiGsDQHroJTed6Wrt0+knMXKd/UFpcXDDjAm88cW9UXAbWKnKYkmYfwuBU9OE5
ozq+k49ES6E1Vz514ua3d5SCq9Uo/y6rCLXvQMbDGqCkHNGRwy1hyS6BhjNVmrN8
uatxEN04KC5SvoTLnvUVPDwJgrv1S0mL35COWgu6wA+Rj7QH577Res+KtwiMWl2k
7xNajBK9YeFz+jZyZk0xsPMdRx0RbAkNuvUqXVPq3GhLj16iB1Od+K91D52uwAS2
IE5qG9j6cJdBGUtb3hHGQKgOXcNeHouI8Zp+VPzZuDH80MQ0tgcjFHyqsc2pw5GW
KZxg7AaIV8sx7qrvgJGfquMuUwwccoCvDRAHyVGjpb8RhTkgL7QdMcK639YyGVqd
vdALp1CTqL5G6AFTgg1FZ5SIu5zzm5doGQeIZbgEQq9OMq9i9g/i+rIfj4uTsNDt
ZuSvqdcwijfOhAQqXcmGbGH40LX82Yu/gUCg3msPvJ4o3tKDbdbjhwytwat5AVZz
6Eo99SWi/aBCRRAbcZX6rm6VFNgKVLTWYyfwFv+mXry++6gz6RXjQAssdqvbMg86
VoxCca/wI1c0lIdIj+el/7bPLahghskOX6595APHiRCvo0s5CGgmM04ZvomrufnS
0Vu782T0i8ofb2XBdEselXmk/QUORMQa4abdecYxZSEtbs+rm5iepE+o+/NtBwMc
z7tWtlbbVrBXrNp4zHGuaP8ktiYHZd3kr5oVerRbxuiJF1SxkwfWqrebdpNOi2DP
tu3gQun3fUrlqABRAYNz0yFvi1FAYccD5By4Hh60QP/qc1Y46z+8fcx6ENajiJAF
fJs0RjR3KxraZ4KJ6H7AJOG/6oPG8ZPpD0trRYb+4vb1j8oLZCCHTt3gX2ymGtkD
tJ++inqLJzVnriHBzlcNwxu6o4nbqRkVElZcHbr3aLNmrEQImWSu4++5nyp8zWGl
yw6JOderHidhj2cM8JXN1Wo2Hz+yITYDyuYlZ3JA5hxH967k7NORG93z+6HKR3ym
lujXJ6x6vQ6zWiVPNr+NG7Qby66vE+KWb8JmYMM6qV/eHdkgTLRka0BWDL2zQhYy
W26mSfRHx3MFVnrrCN6N7lGw5/6dqKCy6IGxIpLfDY9sXttIWYvrTM7IyTGLujei
exq3qaXtShEMfyuDGS8TjvikASRzwvwC7SfMe0ZM7zkmnEk0tkTZa9/GenGvT5Y9
TZmU4JiqlxSXsUkrkIL+aiiXd/pMaTTg+6YvxNpLvSe683nprV/nNYabnuRCoHFc
JWePFs3wsW4Zu5/uN0nZMGLmmTfhPXt2/l3P3SxPtKlXMDrFWmOxddUOltDU+BPW
2MOJYTrzL1hhLkVudXcBaYAE1FP4ly/XXT6dd6dY89XCbfgGoms8PpgNKXgO5UKl
YdKTY6NGdyhCo6BPiksx7iiHx85dT+59BQwrqxQjhU3KLdLj0JlzwxrpakvtEapS
7WhzLmEBMAJu/oHO5KOgCJ9MVu3YMVUdKHgTJWdMZ786qjriVAFYqDsrXuFBHx5j
WaXkXqTejiJeaDGraPLRG70Bcj+IQXVm9xe4XkQqgp/IsOn/tmXdKxgcA6pASzEm
9JPdVsG4aknu8Ib+Big1cgKwSJse4tB78bpCOlOFlSMXxMr6fkUFoD+zbWIRNfaw
zzlquA6/lwFoJZzs2YIwg8WT+o/fMK+Vhyp0Z4csJGgFZG6IPFtOi+AS/RmL66OJ
XsiPbeZBdlT1HtMi8HYdXd/pRcRFihgJdbbhlLNPrGTEV4uhMtwulMqi5Jim8U22
Z/0nzq/RBcAhVAvvLwlSynWKOiQzCnTfpmwT8Y4azwbU3ZZoqWLGBDcxndTfUS8r
I0WLmAKV24VuZWBQNM922Y/9mUMpIshSPdwV4i+ytt3BM0cpoNnQfORMUuKN1Pwh
fGcEQekcTvWAk2rXbGFlHXpG0gGSfHp4/HpsIMUG04vZpmvFPxehXc0vb+nJUAmd
eyyRiErmkV0IfZN9ENQiDbb1Naf/ro3XYfNkPNJCTf5Rcifgc33dXYBdHdXNbnqH
Yjw4iEbHy+E4mmuydsttIJ9WwMYwjOGFwNoG6+kdgYuYgOL9VU2dcvaIp25Z3Ffd
eyENTTEe7qHuJqLMk753KgNA2U6w3u/NaegcyD13XrmKTX5MOSIQ75JIzpGYaCzK
w6TqRIQhdr1mXttx+ZSqtTRcO860hoRUc8Ze//97u68fZAN6/82SfrLsae36KC3P
UXYZH4bbhWzIgok0B1L24z+S3W0D0rbEv7/iaaioZ4sDTaHl5Ct5E+/uaus2Jkxv
4uRPVzW2PqydweuASbExMtWcLgHNYN6ya6owuycOYDQ8wClfIovgXh3rK47u4m2f
0SN4C1+DEPce6UeZIVYInddW+9doRpk7ata0D2wT0L2bbckZDCwvKJKAoQWTr2ir
S7i18HVJlkXR2qd6brxx/mt9cgdtdm1wLwTSROTzoBXtxAYILxZ9pxVnXmLLADLZ
S9inSTbL9RMB092/Da0Tmmzy0Vsp7X0L0KUR0ktdOyyTpTYekt0pORDnJoUmyq5k
skjaFUrJdvcrHUfVMSITTod7dG7sNq1Mk+unChPmUOkjPVISWfELYc6WtrO8XfZ5
OAUzdnBMS1hI8aDfGotomnkL6KX0ED/ZlKbUCxU+3K5r7mEqAiJQALQJhCAxh2rQ
GkEWXGZecKMkSmnrIEpdL5ArSFTi1U1w7odmqKwD+K5PqPm4Z1HxkwBFbX6BZxww
lXurK6fWP3vz1ZsujtC+/ageK3IMRR4uqnkAc1L4SQ9Kv3fBQydRbP648DvuuIHY
gUyU7CisVpSx48qlzk23olcSJncQtfBBoX+OpcepAm6RLDJkctEP9cIDMWqf3KWT
Mh1cs7ZbkA2K5EeXWehsDC+G7jwdDIBPdoxMG2/NQQ5ahLk1dd2GbtfjlBOaimPM
qLM0ZMJrr4Fl5VS3ZDNxnqMF+kjEle8GxPdtQyGjWPS4quTFNbAN0WAFsibQMwRm
Qm5POLHSkcEnI0mM30KM8AYUnh4A1CQxc4ZW0GBQKzHuX/ly62FZGYUakSe7Nux2
B0nvxiCHfww18OONqSYuKcfwsuJx7awxu/pphSb1fhSYlJkGN2mFnm5yGPsf5nwX
7EdUQJCTMrtJdzZBvCdsguPonBoMv1970OiNSpJc3icYnMXUiDFHdwOFNx8XlrTG
tW+SaL4PHNdgmCHoawPR3PcH3tDIM2BNAbuzpdStdtj23PGuEPRp10VOzIkzqabP
eubD1H1uL4RjMMHByEcjvbgDFRWKrsVr8yZzgGIFyP1LT2OCrJC3TYMLs4+FkNzb
oUYtmJNSvkog2meXoP5UhGkX7+wQ0aSrHNsGnVFd4WJPtVW+WigG4jqX19MVf6dD
HvVEDtCUVhHdZv/soYp3alROhHmxAIuwFWs6oU2yQ9Z8OMec+zh5FqVKoj9yhsZa
B+LerKN5mwQgb19uQMtzT8/Gwg56tZJneiCuGaE641y0LMI1Qaoc8MCJYdyj7+Y+
lcEyEuZNi0upH1Ff6VozpNpUWdyOwJZwUNASU1Q2VtNgvFOp+iENek9YC46yVfSg
SBi+zpWcjrR2XyOKqWDaq3P2PN7jV4CvK+wDwtqcso47ZJXssyyk1p6RY9dlDahQ
alJcsgB7I70feTyFQC3z1vdb66aSTkI4pzLUdVB+WJ/8hKOOMWPerdqs1J2Aa5TC
vtWzf3VUn/zkrcicLOvN7ve/iVZV0ddtu+qY7s0wr6TBWWl0IiMXM4+v9s8XeM0/
lZyLFLbgcaJ+y8BKR6rmDzHPYcPtGmn93bbYOxTFbuMSxSO/WM1/jUCm8OMThXii
mKKMPihToiKRc/xfTLLYnmhw76xQTmqyaHGB1eDZC6kC9mw/NMrJZsuXz+rgTCcm
UoUFKWj+FOkoaBvfZ+Kq8WhHGFLbFF8ThhcZgrTUhSiy8xSVm2xCwUvweQzgI9cR
ngBLPYSs8O+d1dgzMAESo8NNA2yCtV2tP0Md+ZM1VCKPgcfiSpYcezOg9mJrgcRE
sr+9oXuyN0Ynuo44bRcdcWujgSLqir7aEZbPwHpLN5UceTem+SCNqW9OxZEhD1Ou
igSHvsICnf3++N8vvbwLcE0PN+Qv9XKte4I+8+jEdtneCjhPsjIsakGMUdoxCWiK
8sz5jUIRkBB66LWX5g6IwAiMk8xTBMccvvz15d0f6pM6u5L+yPLidgFF0zByzYYN
PCz6IpDFSC03L1/gTLfR/St+92SciF71wEBa4ZRVtOyPNuh6DT2VDTOR+1Fn99et
TLsRnjQdcUP8cfoo6clcHHS7kEjtjUYcpKPGLkX7saztcBJ74eQBVbDpNxIXZX8K
Q08DE6p2Cbmsun8yNsE4THBhO5POZ67Kzj7QLIfQEV5MTAvMD3ByZ+Sabf0fqiLE
GyXfDNx9FDau/ap8l6wO9Gr4fRevRplqSobgfPiaSQtEBAlKkg+ci47iKI3fKjS5
BqGSs8reb1jmiiL5hoF2ewoWcOCP9xKbLGEhwPunI7bycynpCJQsJYj7vsx6s/+H
NsIY4TrOApjDKmAcFGm+X+MaPF+diPf8wBYlL0Alc/OYbPUzbo2byyyZ6LR4f/ik
GJ2H2PrT4ObJsvvPINNt7hvYuJvoOhons9KcTv8iFxPmfgaUfr1jWnQb213EPS7i
8mK1PwpdUxd5xRdfTudmhYaAJUMi/DzAlqqVBzG9KZHVPEyKS55rCubwk5SpsZg2
HvNKji7PGurHJ3ItLkwldbzKIL0j9JcirLvTH/bxYelisulKD5JNfzcU5BUCcYoM
58lbkyKBLjsGTFswLMG+bCN4qs3EnexCTqb/CO/P4JAQcDvkGQRID4aJboEuGojI
CeWdDGmK+Ikdf7XsdxtZ5v1+KaU4u7dweb6eil6yYr0GcxsLuBHpl2f9YQYksSq5
yUTnekaTY6lcgeZhbFBn2XE9frSYBU+JnndtuOQeQu6wPNCZ2+Gc3j+S0M4JkeSs
WWlhPXHb8YcBw4tvgTf6ACbgTxPcImA3T720TmDRYNLccW44nl52jC4nydeqtv/l
PgqVBFjhJ86rGcfkMOGmO6Pw0qVdJr6HEM9q5rJXt6KYcRYwRfw+PjVOnvFWwBFR
V1MQJG7xvDJODhRG0hY36Ny93hapeye7C8wg+g8ILRsa48KOLt97N84sRYk/hp8d
MNQx2jZbM42fPNorsp/CRcutNky0NfD5BMKDXqpJWs4tSuYNTSOCFXKlM/5v59RV
MzIRgvPiVw/uj+zRtjsiLu2/D1rzspD9dWWgELKlVRL7Il1tUZqaKWgLR218vZhs
Q4a42kfi18H0+7dOBerVgJxF5WwNOtW1OikNx9Mh42lzHTbSZAQRlSyXuOyHRVpK
A9qKinNlN8hTFq4GtkJHCZSwSbtVw7IqVuNFuKG85rY/nRqfvgBndM1fSes2ZuLI
hgsze6j62tZgJoPOcwu0UbCfAv4gSWpP7VrrAFXHasqsBoU6yXfvXCyAlnHHXmp6
Ww2UingAp0ub69Wub/4g4PCZmb4wEzme8uMQU9v2hsyfys+tgdlrWzpiBwtZ4OtQ
oLtS4vtcsIMA2pxaLjugKDziuuJw58ZC/5SwGL6X6PafEzDjYK3tGrrXMg8GWwMf
7LurRBxnPk0VUe/xSogef9Zp76+3SlSymtxGBijt2Cvy7yh3fAxDRH0Eg0XwMnuO
Cbmb/WijWhfMfBpZxMowm82GmexGccS8UKCfGTq0OUxmaILvVjgP1imialRHk/rd
ScitSBC1OepSZFM00JkHmlCXpFDX3GrUSw6e/dHcdkhrlty7j6jrKGf9tduDD13x
cL19W/HZrQPKwR49BCGco/U4OOuchlfGnqJeDFSMtpjv9GrGYT9qP/O3JubvlIFQ
a/X4CiSH2Bx8urd3YhjkhJAI1zFmkrb/JVqW4Zibv2Aoob5RNUOlV5Qdb5ub1FNn
pmnQhru0K7PHZsz0CtTbJep4A0eerS6ar3KwAzuLdRLyoOSrkdtfRF2NLAQymqys
2GAXj5KOfmp7I7zZ5j20DaOMWXLjn9ZwFhkP7IkBXsGUgS3qmcLMXS5NjVwGliVv
+8gaGKMPv7q0wMi2draWzCTV5VGXNdKqINBygXdj3sxWZXblC3imD4wivNv4u4Dq
Iqjz/H5f9I51yqaZad9TgiaEA/IrRAlLlBjJ9l8FhaXahmgeWc1aQNwYqHgZnkEb
DjdUCZsn+cqOZhu1tqUy98JDlzqQKaFay6Lu1QPkkE3MoTEXdG+37RdqRbTk2ilb
0clGv9+Cl0XU0CzTrtcp6s/fHyJ1k3L2CTw2FxDrd/GkI6i5Luyj0TWPR0nCFV3g
g7AfOeNcEwcZ+YBCoaMzA9RUJQl4uXekSVUAjGsylvwIjNuly1IjNLiTI3ctsJWr
tYocyUPQOhLwKj0kcoOLqC7rRJhc714egaUpG9/LUSA4GhGUf7bXqj0Y8A/TgCIu
ZKUxTEl7WAmmZj3ZWj+LYjdrKkuOg0UjuzoLnZfanVuhpWUnDOve9N//RCaWewCG
6UUnm3+NMCKfgbYE6pqSAHjhSxQPUxHRcgjOQByY/qbSVlYlU+V9Z+s5tsnIlFwI
BQIZOYEDDN3X3gEl6kUwxQBVT9WjeRNe2hPbrB6NU+RTBxVBbLqRyZr/9p50FlhH
wGsP58AietR+/dZvKZcSPsbWIpsfwj1WVn/l02Ty+q6QcOOEZU/WlqjZvehILqF2
6K8Q79tnlceEYS7BVPtX03YawWnsha4Jbr1fM1dt0fl+FWHF+6CBbfp6jgpRgMwK
FKPjPPExb1Zzyr59f8DbCNqzikkRhSDUFhKlncdAA2eIZAxkiK1EFCFVbNwEx3p1
xL4lmZsx4nRCZjxlAIKjixa544shJ6d7XSLiO8vFkJ/RQoHqv7SuQfdlgPRzJR/7
35Zcb3VSCwUMWSRZrEasvocSxtQlOJbZyL2T2/cwsG+YlyEjWLOWcVmu746BTdnh
OrxhpGia0v9g8unhX8yg/fRirb0o3VEwO6MrFjvUnMzDPArlqdfDzKcqHn5Cnxtm
eLiDa9jcd2IERwxubovlCG5J30YDYeqR7Y3EypYcUlOBOdP+NCFlFuTJEumbLMYW
i6hyuQBZNnDdkATDdAunvWKH+H5UMx9yQiyOMF0Jsuu0AURZeCmazQneNUNm3+Dz
VzCDyER1KbHPEXDVfpQzTULVa17jP3eKjKr2tbKB9vDOMdAAGQe6wU1i6nuB9jEj
4NCq5QuazuOQhKEI7dHdsNDtzdl32pQTbdWGHDqm7CCtSIb6NozQPQGrMbcXCgdu
smRJPTNEX7M9YM54C2Pt/qMoHl2ApKv+ooJIGVSsHk+5K/YW8IpISXCX1FQUzfMa
MaxbPwUQWVZEYg2zxqqvXBZsvnL+4LO5QbijauNhg/tnTLgqQzjbTWT2PSpm6NZn
ynV7ry4jdiCeBERzOKIjxvNMZzcykmieHMJ5ldwXrPoPqPZF6MJV05TeL1tNl8Gi
WS3x5m4zV20kPNBhTC8vWCx0aW4H28nRixuN9/FO2qF6dXE9QyHoThJXtII21FG1
igALA3i7xaRBOfutfWY1RqWrj715rN+s4YGS0IJS4UKpfX4gNbT/guu7rU43vzIY
cgpHpVCxVALyGzxBQhHxn8gbqgmEZ2gDwrWIyTQZpr5QgnCo9flrO9a3k24QxwtG
d5AmqYjGt//l9x7rbhz/T3kpm6GnKMeS0dw6idV9SWxSsdyBgSoUxszgkjR5U22+
1mlsL2DPAu2FAiL3wGC06qHBDVYifV8CGHMPVcERHxApzXj8MW5DQ2LF6oj7moJg
srpKc42SFFY9gaqRqVX8ETkxBZ4zWnb/dHH5AcSH4wPyvUIk3zPctT1+u+qx5CdP
uuA/2L9dlj7toqN+AOVP2o3ZFZymT1q3oqpDeWlVNSbgY6QjLBMuioDtxhkM91J9
AOXZuhANjD6pbcWrXRKYBA2DbJyjbRs7lZ8kJWdLw+kB8r0V1KaDkzzkZuLAfypU
G96wwkZimcqsNsD4Oxhdlwxzw59hOmYbK8UHUz7iXEMAbEJIPgIavb9uvbrm+C/e
xnFVsumETiX1jvtsPHGsUiPW8Fy4uNagbXJj7S5LpJe1BWA1k5XQJ4lEvUXUpk+k
WU4Nm9Gjd/JJlA3k85UHm/qD+QE9U8C31LyIoDj+Qk3vcuLiQQ6AzJQC2nt+0TZk
MlFidAELmDaOVOLpkLv0pkpsiAZS7y75LI93pdG/Bw3DABqoCGIxYVY2sLS0X7aT
ic2aUm2wNtkSV21ZrPgp1iKMxQuge+ZWZQVgmw7B9pk1pC1RPZpMjL2jn9xfmgN+
IB4RdZySUEH+mAyv1lh/ValGEUCiSLYRF/Z/+mbm04nFxAtNIww+Zw/xAXV84aF+
QPziDQHFBpkhuo2yvNrxkjg2f8fc8Ca2nVWynzlwe3yzPLcdFsvqqV/qEVczLXFM
rIiIBvgApfIvTirS6qqF475LMTgpmmlq1ssOas4wSf3xpzEEZzuK0oPr8LjOalMR
iexPqWUnzQv35VnNpFmWYnRUexBbPhuM0Vbximx3eqjLw5XfJpnrdFsWpvTPHSS7
S7rfA/grNT+kIYT76g85JcU3b6HlL91BejLpnMDR6ImEgknfmfGT8HJoipsi3A/V
PVGqKrdIS2jMsm0P0AaJqhepSR/KPgP1QwriAd1gOhDTyWUHQ9f2/tlA6EGCJirW
uCRkxK2C8R4xREa3ApmdiClPGgGdM+Bz5HQ01W1seslgadKtARB0Duio8E6q2EXq
2AfnW7HvhnUdiwDrWhVDt73N1AqYxeUwc+jX1+5LG1h5Yhz/fMnKq8qeEwnnP5QB
PjajsLOuuUJvooKX/1eoHUcNoya7vbKc/NlirlhfAkuKCBJmDmsN+4IeB9f2sHQ/
2REpwCzOLp3OyEboF3pNCtGvVgLDOfwHuj8Ac+1XcmNJ5PWESLwTZIPi30AU6m1C
S3XXH9W217rHXoeb82m1NOgn8+jrJADOjFV17vv5v1tJ2cPZ4wuKUQe8GY6VSCCY
cPSgbQ9p6mPmQnkq1vRqXQGxWGfgxXVYrL5NLI+vsGmWdLjJ0Ro8hXHw2SgE7Sm+
Ttv90nEt8QmQEjq5tjp6R+C8DtV+pMGr6x+E4cQEO7+BIvbqz8spPQEOI7x2b3b7
B2qhSaamI4pIFp4NWXLndge/evaw2ISZLTYl9lEAQH7zGYTvlsye9TeiWwUnHndu
DVtxEJ/OuBIOMOdyhqYFA6q2Da8T/KAxgRFIOhbtXmNFPp9X1BNwQHOhjML9t9YC
7UIbfi943hHWerFJup1Qg9eYbikfdtSuxFSYSahQmf239jQnb8ioIt43fsFnES++
cw/JEIgAN0TvRt3zNBK8AimbodcysjJKyzLQd5f7zPHLZ7iuVDWElt0tNeJyzfyf
vnyoNFJ9gurGQZqJ0/N9Ue60NT2Jodnrr/bzI4ZoztKlk50mChK1jDa4O/SlKSqO
4UbfEAjj9pAnvBW9QnpO9BJ1QBwdFSsrMRD2zMwvf3PSKz7jMV1SG6LbRbf32tY3
dFlfUk82rlCk3D3I+lvchlLHogd7ms+lpB4R7ggAI9+4aj8RYkVo13LYxsfzuODr
1zr+pKXKj26xM/Dquq13ecbu62zasyMJaO/KbWox1AR7JtOW+ZON6Mr6E121XD3G
Ak2ejJOEu/hIkZaNJpc7xOFBemHC3o3g/Lhdqg5k8jB5O4oQHxlfMWtPY2d0na0l
HUC13W2y63gSzr5bij4+73VyUmEbS2thmTZDCaqtI0005Yb4MsHoKW2mMw9Puaxp
cLku2hDteYcWCGdSnHwgD6hPOzEpsIGSHY9NuEC9OhKSJjd0SFk7kYPtNCVaE12g
k1aYHIMvOirJBEG9UEeO8QUSz5QKeneeq0cdHLwxt3z3T9OXfLeH/3DHwP6xdhTi
YTJuSvk8Xltk1FOqUy61NIVam2qZQ/FvpppYbLY3mSgtsidPGSXYVSf2XIUhW1UD
/Y1ts5DUNl+Lpr/GdwvnleQ56TiZzGEY4Hg/GatpeNpy3LRf16HL7JV7sXXjTlyf
XxH2F3phakooOHZIy0tuYvc36+mSQY+fknmi/1KS3UZf7nSqWJYKnweUNEi8iIFk
KAC21WW5OHIpaieeIuRlp5VoeXBa1NZtBvwqKyri/hGg/YCIKn9nDhFCMQufJVoN
C/H5lAVA5v8j6Ho/k4l2vlmxIBdGn2/6Y4jOL9Xr2FIerqIvd9+xXr1Kt7lzQcxZ
f0mnQCvPMEgt7caujsfC03uCxs1IzEg140UgEZ18ukUfD4+4f5Sk9PT8paobk1qK
ZQR4FQLi5xexYQIkCgiKhPr2IsqLJocuXBJIZg6t9F4duqz7fp/QslZ7gcGkZpVa
LYV+CuUz0ii/LEYSGLkX1IfI65ZHF/7iqYHP/+sgIHCexZCY+043MkqOLem+gWmc
2X5rf6snh8YAemXttzbbkHYwAy2bN33cyYsppAQv+RVRwgdOLQxuBd/8GIvmH96i
Dd2P6r/iSq7m0ieguBet1KE7ZAFsrD/myjaAJlDFubSAcRE3O0peRaPyM+q6lhWN
aIBGWu9M5k4f/aUckoU/LVSf8OE70iOk6r7WNUBvVxT4zZmpFHM1Sr2kphBaEfOP
1nC1Ky6KpSf+/yd4ST4AYvBAqhuL3dF2xSsR7k4wLLcr+4cGiqmBHdKrLqyXWxIg
EiRtQOY7QMuy5Fp6HnuUpDT/OHYvzYqCFwyK9BSIpWXraJwxLhzeTF1MlTarN/JD
33eknbNFdpVCEaOA/Jv70eiQFQJZwUo4GTOq3rWT+32PVMsyW/8i5ZIJd6yVLB+a
y3LKqZHlyynEdH7Z7Zci0liFPU0/8wvsB4wiujAVxOua9nBFNHp4HYbQAs2yuWHL
HEUWFtYPQOd+TV52UTyWEFRbxwOw7Sl4Fo0issA9gJhqq7FKgrUyDgbYjVnbjmA7
ZRXjAI5Jgwhjh4Qzb+54CVQ/TPnN14T4X76H4PQwE29vs7GGjQIU0O0TLCCJmycc
zySfsCQjnRFSrDQsutA/unGwF750eG9/gJ2q4rGBJUqySMe28rDqReGh3WUMUHCY
aKwsNp3QqiEVesMwJwa42h8wDPEELefXj4V4w62j7Qy4meNAVHH331sR1FKxtqjg
yKzKhKwRzKLsbxbHPF5LtQv/w1UBVjyYqGJllYo0IkTHnoEmI2yzqTzidDspL6xw
kuYAW+LhisX8RIPIohml9E9cpEU713cr99G6PidPK2WFHgML6ygJvFdzhMd8jsIi
OVzdtARZXmBluv7/AG3ZVqy+xT0nVIvfx5vFPw4q/lFpWGK4kb/V6peMLj8IHIJV
CCFKsOMHp8mfEPQshVVIRAkIdQMa6fWidjw9GYjYGq6LT8DpGqfkSAb1ZbrlP/NW
cRYwGIGAgrjqHZcHRr3sfjbKv84B2FZWXaQMN0PYSLy5IFW0JSrCDyIFII1Hk6n3
4vxUfH1fEfePVGIm25vu/QydarBthiZZ+Pm1xCbztPHKb8eE2UHviHtkznaFCeLv
IiD38tgJTfkRVoJ9LN9jz1+LpG+dGDgvNi5zroMtTujQm+pon5Bm3VS5fFiQAWJI
MLVa91vv3rEUstaSoRD9VNv+g3ZCWy685EIXzqqIa680gOmf4WfD+B0O8DTMYA5M
olYKjOcrvLMEoZXmISYX+kAFttzrkaGr5i/l0mcZhaPXn4IzV4Mhu0L48z9cRRWb
Du6xxFbzK/5ee9uUwVqWvDZ7i+CLKc4iknfxY1bOkVjH/ccHJMmeC197KgnSRsA8
yAAlHiSvi0mRMaSprq1Fx+XShH1pwUjzI/V/+spyXVLGvaTjqM8mJLq8UBioM5Sq
JiGrkB5+cW0XbIT6N7yvHfIIhUpm0VCX00NlSbwBBPNOU1DSb5iNPRsba5zGuwxH
hmxj0ivgxWwb3lDis4VOBlJk2rO4slKb0VgfVOUhbl37Mee3TfXbqVKdg/3F4Zju
Cr9sjj6Jq2ehyRbiDZk3itTp0V2or4Tf6gF+1lblAE0Ptd7oAzaZIB3PE9fndiwj
r/Wh8jBnyHe+AfG08jWLfE2LZ6SFSqwZhnIgzzQzDEKEYhz6P5Ei16GE8mDtZoSl
6TECNiW1QOE97nSMIGm3ClShlQZBQ5+rMBotSP4Tat/c0Dw3N+n0L+cqLGNMjt4k
Mp0f8Wr5SRCCDNgBlk1O9E1X6n7j5VnXY8l591INLvLotjNDOyqvky1oUeDOva+V
AHwziW9BGAAMSKIMUKJEItg3HWaFp+4p/Oy2pGs1m39QVwsOCWv9r5FfUlE3J7cb
X6tP+uqNVbrkYVI2Psjrf9BUI4NoXAnH1xFD5svfgU1NXVWi4qdvNTkIV1TALRI8
pJdtIovSTDWw6XK4en7qyL8n3a/KlntLV+8xyBGdhNYAWbf2JH6+uFmhUwC5J06t
6y5FW0Zv20brEK/J2yHkuie8yzvE6R0Ld4m3T6VCPx7+0CcOMELGcpPToINT/1LE
gqAU3RBIljSO5AUzClhLoiLnVjuOQrRrrYg1OxPWwnV/ZXuPv/7I0f5NCDjePxYX
eDGOcB2/rYs188i3qMMqwMvN+J3dCXVuSgMLiZoS9k46s8ZWnMKTVRFxoNcVxnOH
rK8yIsgzXPrnAhbex0UR70uUyHbDkU5030pAdLJe+KAt7haTTqwEHvBg+dQk9Eq0
F/UCkFNe5bceSnshzKra7o2ZCtolWh3XxcYh47i9aYnTwxBw2+cJP/H54MB+cmOX
El0NqmKUax1ECiC+04mG9MwJWnd469oxwROsOX+prtG3FqTLqRdqqEqxAwOeEuEx
E+8akDSsxL4sOBS+uX/IhBLA2zWR5V8iptUt7RfwI5lAlngHKVHc7r7GUDVK/K+T
SL1hnq+Cf2xbjGkyOt3NIQuo6BQ5STsUfsHm+zgrhVf4ijWfT77KRDusvEoAfxUC
PdOnEcxtiuVJ8OccjZeBG7oBN/fMmNOchCRNE5t+YfBMDc3/1FhypHJlfku3YEG2
hJUHl7Ly5lM6YglWlff7L4+i0DsuVmYTYNbnBLX5rrU9dyq4O0g5U+0jIjExVn+N
/qxUwsX4dfrjno8sCu1tfQfcIzLGe4XfkCXtGqAQVVm42PvUHbkhYyqCp5Zovey4
WlXYOVqVz/aoj6gL7STX7TNPsUM9KQwkH8aiI50mtJv5qFGrbeYmmUbpj4jSI/qt
uu7HMnk3JVA0QydQk5VQEynsUYYKQa22++92dn1UIkuoFBZqegTavPsbmLaNdItn
dIMRkx6TH+r9AB1Hb9wCYQdI0ZL0/09uO2iHolkCDg5+qfCf9aVncB4mUZFuMeOZ
2VEVXICU0+NEPIT9F6/RLTEhxSQYHl8a7G6AgFs4b8HAm6sYURPAPf/JzgXiyuvA
xoGGy99B3ru114GwNGLJvOC7YhR46u/1wjGTEnHvXYNcueb6CTwgpDD0rv9WAW+B
7BuuOtZUDnyq7DKJnXQbhvDfyArOjkN3hdlwWKSNTZrEhMbgU0n4MWAL5OwOcP/u
lzAEqn0+jywYOmNVu1gtpHRrpzj5DDPY5PaJi8Vu/V1ZjRTOPwK/CUwTq9g/FaVO
uzKSB5xCqcoyc1dtbmFUCxOH1L73S+1wledL3EqdbVg6APMEEXGhmWFXtk3uw0sy
2w5SoAGdmkBGfNI4KIsBCbi8cjKOrKBKKISMbntDW1eteP/962AHDNDeoR3xNxl/
MlrCPSRgYGKmUS/JUCcHtF+KEHxYF5CRU1/DrJXwrt1UuX/ZmfNq7hKoLbP9zSVO
+Nm7+L3RhN0nt1JeTNzmqHVz+y/umtgKv9SYbMESzTDCbRKjrxNxK8pEs3qw2+UR
C5wAjhe4n6ye7E+dKfB1/FYOuETw9rnKCfwsOFNE47wNPFX7EteGAgqCD6zrXLAL
vHhPPm4NEuFdGyD3ud5wnUgOBgejhAgN0MVlnb1In7S2uINcLmIktNCkI3W7IbL9
o+MM8oufrQmx5s5Fs1UBbHiilGPXhJijnd82VHRWTq+YCF95RHhian4BLr/C12p2
CnDkCMrGu7padyr9uhX+qCl0RTypLXMqifhv6WKEk1YgypRdIvr6bdykiNbRtE5z
KJEw1RK0e59zPd8/M35xaJopQZ07w+6ryMVx1gEg1zjKH6BvRSMm57wGAg4WNw0W
ag9+8FBJRX65o+UMbeFyJFGK7aJ2nPhIgldiWeyiwzf2eZJnir3vdUdL2zDzsBYG
9HyyXGpZgFylfflFVDwEgszJp5tSY1NR6uwMN00P8exHsNSQ4Y9tL/d4g+IaR8Lr
KdIlROioP4pjA0xcdLged/ythUNRFUOTS+Stikd+7QbRR65IM8f6CqWlKb8w3tK3
uc7F8MXBBcitf/xYHA6Y7LrBcFM8NderAxRLsLzDT21PlzlTiLqmV44H5dpq++Az
sdZSU1gaOsOCJGxMJSxHcFyvQeD7cIkGdrxNfClDps09SuHR5Gv8pKPyhwwr2qqJ
+NTmaI1yc0whf3XZcY5NTpmA3BLl32R0Mb15gFFbemWAGnFARwApixZ9XnGZRoSt
1jLtuZ3fUtoEO7bwt9pv+3hTEOqPjkqLiL181ysoQmSeYY0LrieQqcrjGth/4GG9
PDfPA2S8LckKmvx/DvIDQlFaw6eyoSw1p1guBEzOteF4I95iNIqMxJA3KPa/k292
be/LbnakJaPPrBhakOJaMrvc6wdP07mqNT5/EvyYBAAXWXaKtSXRmPM0JHzmO2kY
ZLovw8thz05J0TtDS/G9WOVPPK1NMLoDPjrE5StX9goZ8FpuVJlvSDjMwWW+E237
m+JNClAzX1ed2juwFMzyy/nFbPq7eSwhyJRTKQ9JyixTPZ4YqsYIXBYLVxmSpn8g
GUJgX5VLDicikcvoOpSjBeF2Mr9NL2+m1OKSTGl2FTTne+yuTh589n4Z5KcrLKR0
/5ekl+dI8Ws66KpXUet421fTWUYwiUrJAQAuxyzLCM1lQSLQ8euiXDQ59SVkVwF0
8hCgbMWpGQcEFYLlhgQzK7GvzUDWVYJkW58JdodKD/Fg0LSA51yJ5hknI5LYCAxW
iYH4CoKrNhJUqQmS6ajgaUbqqQAqLPLEjpiY6y27jrTBVOSmkec0L7Nu9gj9jofJ
PN9G7l2ayYeZZlZr5RcSPmIb3g/hmmghW74pkDa+CkcqBjHz10YJZL48u5BEE2bs
KbSBIrjw8naT7gB8HT2GIFuLOgrqcW0XwZXmCs4suzDRHmd4a5M7QWDwrZ9vN4GR
Geeia9LXv9QfxNceS7L12RW9d3dP5aPGJt9Fcy7zzfS3wrwN4adbuCcAsnDSu/GA
QYrx1Q6L5fUHcBF0U68eD8nsh3kAmFbnjA6sNAHM2fqoxYjCcCpSDTMzug6MBK9G
QEBxKIPUqShre62+8AOxspGOWP9Hat/V53wALG7NbWB15OlkMRSMPAbuzGAoTAhF
NEemVTSCRiANQtFX4Qn9oq98odOwo7dftRJ3fRHlASprjYDqp2s2pMhGz0ztacH9
wicmecPVf9lTrPJ77pPQD39didoMqfI60O1Ie9Zm71dbBc+r7dG17EOejzRhwW/0
3q8vhc7ZfYiJyxQdk1BQ9q3zMkhYwp/AkyLOSVdIH3gU5ZLv99lSw7G4kOuAzx99
GIKVsjqCGZdt3I2KFFq2k5Kry9xHJzeDsJx8S5y/qt58HSc3/UzqvVuRcAkhfJXi
p/W7LiU3E1lWi9qJYwYNBCsZOeK7HLGBpAVLOQDpkehICyA7I+PD9Jkhah7f3o55
azQ4MSJ0AnPNK0XVmeMzK1BPHX/gO1VJD7rHZTNCdHli9D7XQIsogYGbD56rUT/+
KdndcBlbw5zFSlEHaTeJvEzRjq7V4+Re5gZbVQakf0AYk9ni/WEZtEKJq/bow1hh
XN+Nrc5sm+S6/EnzJemNRINT2Wqa3v1jFICDrn3pojMNkIph+Np4LpkxR7PAjk7L
VauBtzLYGPB/ayyEvDqxGBsbiWitcQCslAJF10a6ODiu5H9oj7hCN6EbyzWyKVrp
jprVgm/FDZhvkNR+yynk/45uTqXecwd3gZ5JYnzEIHKzFJbGCBWmk8q6rflLrchI
ONMWEj+xfgASmFJmkRjE26krJDFTQLMG3+ndpe1GIq/4X+SDHCk5eFvH/9n1mDHP
xIuoz4MGoLl5Bruab6Jf0vNAyzvN/O77GjQYbbPhPTFcYBh/A09C1WVBgcDcFGZ4
vwj1Ga2p6Lu63sPLkmTJ2EQkpBd8ze85IAyJcZfWQXs5SP8pNJUKDhU+gNuOyE2b
YXxScEDEa8zRWkvCYx7SsdjY3Xb5oKYewuISuK1Iyich2pTkQM96l4bnzwyYDTLH
ta3s2u2fwaW1gNhSRSdAtBky4U3NyPTPgpqslNGfBZJ3pfAYPC6mZmJOmEF1xRo2
hmSlW2xD2XfDvo3bpg2KdZknDIg6Mle/b9LZ9pVZc9bxM1zZz9XXokYq4P0r7qyh
gDjanSAYqPmv8967Lu8iQYznm4XOBQM1MxWHJ8gRNBWjneN/8Vk8U3468H6HXJ/7
J2gDow0o/f1kDhrtLyTA9l5U9aPxxUjdopE9Vh78skjc8RYRT/ld4bd+X6ma2ypl
vRTvCiNj0wE9S67zmnraN5m3Oybv7qkGHPlQWyO8+OQJorvoLwb+IxXXADwKdAQA
1B0FnNjzzsskI6kKf1a86hz3SkQeVI6xRNT2Y8zH15NnFhbStD3R0AKUfG0muUNB
Fa2VPCBm9ZNfVk+d7xia/cxLuiSEKWbZoRzXK0UibMEdQyGMRifF3+HcKO5xEOfV
ki552u69K/8oqaIgmZoR6N/yFxEEyRF3skP6phkhbQqBPqX+0aZ6ds2QtJGXG6jo
e8Zi1Bbx0PS2DO57+7T+t9Z4sA2qvBB+ev7xHExlvUjiH6R3K4UTBwzmXZK56sT7
RggKbKInKhOZVUemnCPZU7ETkw9U69FpPfYIypwKD5h++d++Ehwib5jgxgMW4I/B
PUkR4Bi9Xtu8fmDUFp5aDWARcNgTP1RvRJqu30tK2ALcHojGBSUGAUtMDEKfi6Nv
Z9LKfT9GSjvzoE7hRIteoPClwbRJqgPNV85EivwZ6tgpRlEy2wRMBrbOXGpCrxUb
wTSKfeX+cBVbM18JJF63VSQs9Po7QtfFP0JZ2zMUcYtuNSlxXRhWiLM+5XGnuHWP
EthntTefEaLzPPQ5BZ8cZlCwAscDgqsWeSDGNGoYhVrqJuToSNdD6lcuZ0NFG9ug
bmuVsdqGrHH87W3caLWQ16x8VQXT6ODr+FfiWBM0FDciqNInJQ4JH+r6jRYSJ300
bikUdDy9oYsoWrEGly68jxcZfmJqiiKqpDbhg2DgoWsdextYuGhI571FW9fzlWmk
v1tMZbC0+28CNc28jofmF8TNlGTPJYAWS3+wXjvt9jwHhVqPzUc8y6O8AoANt6g6
DEOh23dW/WEQpz8RN+HqL4dXQ+9J3QOKonqDxZXgwIUBQ0X8hkb/esxsyxqp3joY
WAcIGjKqqSj3U4u04yHDCleSwfWI9wkZjimuAr2OlQPoSFWUSU4hIRS4fwsH6RGS
HJJ8EEgKqkMc/l0Sj/aZxPzAXHa3zpKCK9WGJrl7ita0dUTXiowq5VDTLEGCHwxP
rCl4a/iT8QGu8IHn8CFgOETbt7ztB9XEn5t7ReG57KfmuWUMb7c9WsMAGGkVpZdB
tmjd64klCTGIJSeCeIc/ZomBUoFIH3KgTwcj5bR9OH3A5puFFaGfJrTDOuoJboum
TMhhlWbG+XNCUIeXlEwAuvWJXVyWG8/ub7N3A85yjpithWYZAE20knkS8chRCJrQ
6e+efuXrED0DveqsUjzXPea56HnjO8qu/4Uj02096VzJ4eNJ0QBrI/bIfzL9sxIi
JRJjacgn2HEXUttDfF0s2eVCGw1Ng2oGQBFMO1ZR0ajpVQ0nYq2BDTisT00A+0lz
L0P2WJRPv+Y7igQfospDN0ZbUCV1id1lTyiy6giijyto43SYbeM2mn0D8pp4R+d0
fQwm+pK/YKeJiyD5xMw+lx3Y9P1t+0kLTc9/EXCZi8Q0vry0jRdkISWlDVIKux1M
gtSWdpvD4pqabvnnY8ra7pg0qdstCGjurQKQJQ6Ef0HlP+4Zamc2p5JzPWCSJyI6
ODVGovc/DWpI2fxTZIk+pFHxQZN2vQrxhxjVUtQZFY18sikJg7BHaFzSfFYCzjp3
sDeju9dV4/PggtOB8p0/hmjnRYUzVr/PkiMU8qFbQKPhhpvpBXPc8qv3mUb4EkJY
YeX1lFJbXuRH3M0AVVN6Inr2u/fvaJNk47YLJaeddlEJbkAWFNxu3mUc6esKxv43
3J8WxR9S94tex9Z2CDQ7Iw33r5f+DAm6x3KbnIyTAT2rRcGvyy5Q+44JHwZ9J25k
by+tOEKjqaN2rkXNYgLs7vwJWZl3zk5CmiRhjyJHXIN/zPfcYPfQ+6yv6UJTupvX
i/inuRogqfNCuRlBze8HDWk5D3azVbG+16cRUWRYOuR6HbNfhWCdlmf4JywACbx6
FqZGEa+cLhWxuH0WjzAwC89s23VKCdMM8rpNQO3vKMcf3vODmJbozm2L3DpMmhwC
LWyLBYOykqFQDJVoJWseiwKyNCnjL7H0STNBOyFk4/FA34I/0/wJkcyu6CU3LwZX
LBDKEZGoLDg8W+k74+FMf/nCUTKjC/UzZzKW5jMTKiOrect3mMxfbFqCwzo/2and
5vn8c/yaLlOFZdv1XwKM3K5rdqrH5ymV1Qk1pCAfcXEgrSjGAJC407b9GTfqA9qH
BQ9HJIUepwZrj2C2n6Zql3+OcfEi486sGuiktwb8R5L0ZvK919U86aMoo/3LU/mI
tm40G9rebOTv0osBnLLJgfZdQ6vK3XHbQ91wg2Gs8rvgsAW4LwVzU9bc5QnTz1j6
pq2k0ipAx1IMVpy+eYS/cr0PtBwlsqV+RmvWbSI/5BauZihD9Bz/8d6HjPMjAM8x
KKqHJ5Mt9g4w2M2f88ALJhWaIEqiQnnZS7CWkhfEryEl7IiqWRs1RI+wI3v+dalX
L8/qjelnwwBBbsv5n8HgmN1esHoPG8Pb1b2pKB0H57BdsCxg9JLvit4JsjPwQKhA
6jxwdXiCv9SD06RQVh0YU9Hvc31WBfPlBU2TymcpUyzMoM8VkDO2Em7Px822JmcO
UgW3WV4b/qXDdNCMpChUvySVwemCMbBwglZwtdY78NSZb38CEhTVg+UxnODsfg8I
MeQ24tdjwnXENM45+LhPMYBuRe5W687qq3sIobUPAHDvwvV3f7Pv0S/H6C4lZTcN
UYnY8MioG6OxT31zULx8b7td9mTzRSBGInc/NhY9JRZ9Hnd56lqCv9gX2aoS9Rsm
inQd9qXiVRZhmPLrsfJ6wpFq6fIksNchxMFnupBwi6f/y7L+iGnhmcko+wt3kRiY
sIJ9YMseyiXpKtrKz6wfXhZybQlbMZ3FnAR4QagP52NgfxZAokvDASGvB8hJ072U
/rzb8tU2GIT1/Su9X0cC0LnokE1Z7zxHh7WACdPNracCpnK0lu+W9FJorQ26vCPU
WJJJzUsX0C7nZS5WYlp80FvfDNrGemmfsgul9QKugXMi+ZBO64cBpg6tLCVREiLW
D/pWXFBJQ8ppVHH/QHzDefiisrjwbkjnyxrAJPJFAni6xMSrKROlY6Rd/2LDv5lO
YEhd4sJwffzldBa6tOE9AtF92aPAEdp3fG/63mipzohvBnDkXQpUYFRr6ZY4GyxI
sVoA2huyrSQHeTaARiynSQFOqNdtmECa1S3jbPfuil/DP0Qpl02Mcb3Pc8OXXkQt
0MOsMHygwXFyipxBnylyZ1BeHANzjqvCjmOSe85CcNHf70Md/7BtacofG2tLUSHd
ZSMPHo4Hk8hf0W8F4acQ24y/fh2MaGw0Z1e9RUW3NfPOt2GanNcNJAdMTk+y6gf0
gGdIAsV9imEOIConxnwXzdzgbNTtphzrhieTgqikMPoUYqrpzqeKSB0X6QXd9CY8
5pO0o1FFWVPeMomj9FgETX8RlMi3Nmz0rUsUUtNsjBQJTprsijTyNkY9gzMc3AsJ
6WbHyJDWLOtIl4RZ/OAwBT/HtWpznCWWt9+RxYBT7HTjtF/DFT+VcuxnL0l8lgB+
qgzrMGcjzClr6WueLu0NUqqIhbbS3YXZ7+qrpX2c1bRHVZKqhV+dRmjVN+DWOAhv
XYBtczHByvHw77pyFm7WJWuCd3pEGHEZYaIhn4PujhzexzlJvt+wisnByl36Yla8
Fx2ycsd/MRy9G0DdLRhkbse8Rjn8hjyRQMENqQAzbzd3q6jxDrhqzLBXHXDX7lYS
7kUabd/eECDaGNbRcqp7wTd6a8dsA/E/oBl23pC/lwzLRL4Lg5GwpR7wNH7XloJu
S6O9Hl89kQuimZ2b/om+sezIJkuXWoBatPNM86iGib9tV/ytXCypbb+oqMjGl9/g
4/R6i/IDwvIC1gSqnAivBYr4uxkf1O4WL0+NQAydmteirSIEnHcMiZAV3F17/T8t
eUOmRVqfollBDtWakrlWwt4Yb/5zY7M4buHwP3Gch2pLXn1FzkvcjwvCzvGGV4Dm
UnsOwe1GXGIg/+lX0uFzKotHvKFJtrh18tU65QONHYFw7Xvy2gIBjDh0bYKnPdQK
AIs8g72EyfZVL8YKAbXB3nSRwnG8kCapCkjp3qbaUIoneriWe3+8U5mV/WcsCsiJ
p6fAmfJIIQXd6jGFf6XQiMaFd38GthBOpZviqyNkCK13fGy2Vq1vZNSyRCiS2xtw
mkP9g6f1sF0YYUknKG/UneozRTp7OUG9WBWfSeJdqM5o7TBxuafOFWBL4BeyBOyh
oReKohyQKIuSuz794mbd6EHpminZiMHAVQp7RzVoJxp2wG7dI42vTfQkfCaDT4T6
DBykR8V4Rg5zszpF5rci2/wB7fEnYigCIClrE7gMnGXXEremvfziceCPr3FKNmai
87lYukloq2p5oIXjHf/UCc3lH03/20n965g+ENXeeQFmS9eXjD7PEoxsphHs5XyH
eFbQic1sNEkHF45bLHzA/v62uVk0Qns7x/U77+wVbOD0Z1+43nkWWsrEH+SE06PE
IeCbMezziiB5KNEL3lvnue2mET0GwpJcE6CZKqKZGTkW90nEkyfN4kXPtncdDwuI
lJCtvvIZ9iHhqJGNmF0Y6+GCsP1+wQtrcLNqdg2+lfNVwRfXkOIGjZRjs9zAjiEQ
UFs1wbq8qCoVAoXem8o/sBJqXVoIGdcUXUcHDHZfjI/HgmudZj71Tx/UbGoCvKEB
k7Kb4siwMzwnm1QvX2cmKVAwCoCPaUWcVBm5uZbZPEVrFrePSJTUQMISHb9fb3Or
fylkDYJrY97VydpnRwzaUpWXM97UwD6qFEd9SZ5SBqsC8uVTSG4l/WZzz8MQZGwi
r86Kbxn/QSshGffVcqsk9mU4KzoBJGzUojVFueizK0pE+UeAye5Y3fN0++JTJs/y
8la+WjGVxgX77F2RjfJhyHIDxC/UaJBgE4lSdKhcSAmFW0r/Zz8qar9MTVDnZkgj
lhO+DtJPOQ2wReKoOe2X3j6pkLCPdCM8Kf9rEJ9uCZRxXsVWM0bCcjEVjWsM7fL/
hBuygReFbY3PtWM6nq5vjvxL2tzqBIETOgwYUSmQ68YN20isBtRPHsqVgqVMujRs
MFxQ/Vu1KhcJLSjs8OZfkYUbvpololdckSy3vv3dheMWziHuMRSI/KSHPm31niKP
ETW0QNCVc3LOuxpKJdcgmXnkZ9lv5cl3zjmnz/NKvic/1dFLtTFuFvC8RjE4OWhW
gwi5wDolw/nQW5lgPWH5VDF3DUXO5OQKsFC0dQpI53AP+Ox/Kriwkn1Ywydy0up0
hpIqrNq+j59pQhEZj4gggssmLufcdhcECJdyNsR9ZoWKrph3qBEPe2yW+pGta8lM
SMHt0ofglWGjNs90PSzwnwshZWIecufu8hOkuIhwpbk54LedrmONgiRgxzXLhdYK
X0x9O7s+WIwwKe9qYJCNW6f4C9Cz6ETvfAFS5B0f3ElXksd3kDHgyDIZnxNIA3QE
KW1PFk8dYSs+ybHu4/qBqnf2y6zpMVj27Pkqg1ccIhEAjBSweMAAKxBDZJerOd6Y
7indYobBwskXv9ZoYJCEx5it9RmkqWtnqnrAE6sI/XT7iiyjMgjNFH6hJ/rtKEBe
+XlfRFKIxLPGMCxvCt4zpgEWpk43oK15vxNK2zxEzUy9iywRP5bbHOa+MZ5bDEZC
c89z9T9+8pShcoLV1ITi4fn+Fr15NJl4NS9NQ7R77QIyJMd/LXVS893/ShCrb663
IxqUppoDzthT3DIRnPbECjtd79F2FTRFeoqIvw+iVmCQGaovz+ogHFcQ8VrwtvE9
EOcm/2L97ObVbPnevSI5dcnm7dVaR6m6VT27+QsLdMg/LHs1iGJLJT9uiuVL5HcA
qX+I2JEZ7v+XSOYmKS4ghzGR0AG4k2A1eKbQ7AjYFGqqIvLnz67k3z6ri/aWFp8+
ccZjFcsWg/hXniWhnKOB9grBwLyuxSijL6TyJ6xIonvmViZAz7SVg3DM+fH05qW+
JL2en0Z3DmLU5sha2guLdJAKQg4VMeML5CQwCt9Lo0RRfAHmg4n0qgdoxKwlWwYC
oDYJmfMcikNnqQ0cuz5Bo1EX1ojT3U5hj9f6u+cpp8oS8thG0F/393N0IRmCKZTY
APbnHdfjDhqZw0pLCElO8SxYuTd1KVZTh9kJ1UqfQT4ZA2sqxsEorpe8eCjNzRvM
xSvIgTQdwiZxJpsDcrPKQ1jMfkL89UIhhAvpU3JTN50s8aP/QSS7N0ugUSm7rBJh
wEMjaw7Kk91R+cRdAYar+xhc5DXmmATYL/Y0YjDRaZleNrbX55qAS8o058etXnuu
ljBW7/d2Pd+vyF2272GmdjRLg6oNlB4Eotl1TST1H9qjAZzRES6r+D1F1pt7mVk1
3K4XQmBoa+iiovnxrZZn2HUq7v3RGP3/SIGJ8hBD9OTkwENWlfJvkqylVGiLG5Na
7xjHu6dhTtCVrc19h0ZA5uwtLWt0CDN3aQWsrTQyjUCyVWsI8Y2xLQ4eMmFDLh1c
SLOBjaGZP5nsz999nU2lj4ByB2T+FN7/0xBu6dclOT5bOSx4z6oZwqsm7gsSQXIW
+h+aumdOLq7nInbisBP9rfZMAzlilB6AZ6ATi/TxUau0x7LVelqR7I5/wE0clZMO
3zmMj8x7yW96fNOC6QBfXuqVKr5hbf2cWqROoqmVBzY8nYdHFJb11G1rDs0bIuSk
zVyHzea6Kj4PMdONiGqx/AAES3HW+drYwOha/FTNjhjKeig4PXqO8rtqeAy2fx6C
r1xmlViz8c3tiiEO21kHg7PPqy4FROjalTAdtqZ+sBblnyOvB6iKsbEVdGxFd1bN
AkwjIudXfPi2/bQ4thv6qH+rk/1aIMeY5A209+jwUTSTgxuMXbJpJLvGRoLkCUPi
XiI1RUw+fceMRieh7IV9apFyxmAySnS6EAjImANU1oNAGjSkCSqx6qSPPLTtyGGO
wRzGs5xGrXGYcDBcCUhSKAp1S1Z3d/JCOw5uxr7qcDm8JkIsOwghqSgefnqa/R+4
lMRQZygr6lh+NvQTmRvLK/p/2i3yI4P3iGPRL0nW+EeOTJLXYaYVKu+mPfH3AOG9
FZ3P5TS4RLzUKx/Y7jQABkp8n0j/1kaA6LNpSVbus4GERP6p5OmAklA/0lzjlzJt
scDNLnUepUdBMH1q18W+7JWwPT14IDp7A3TmQnO8bqH1NPU+HMb+CBu48FWcxvN3
AQyMLbWJRv77wRCTZqd+vwfe69hAHKCcJ1HRHp+VQLXL0W+DLXAHf3rPRZqV43h+
go1yTn0OktumIhMd/LruDD7dx6qgPTwWYBNwDubyfDaqcZ46gKF0TAEVArem/62v
kHfJdL3Pg3vu8/AzAS/UJTnOkLux2XXXgG/tBg325V9nWRYgss27CfG5gbmmEU7F
djyi1Nb/0XOkqkCNy+7GkHGzBjyfv8MqSVfu3GIof5zx49Jczh2h5QVScrXCVbBr
Px9CesEwv76lPzf0BSPAOYWtjOvgJxdx1KTHOeUq3bD8OKGbvgjMN8l/4+TXUaIG
Fdd3NFD3n+xId7XxbmqTwT7003bmN97GuRoesaUf0W4FsSKrV63SsrMVKX+Ak7wz
mls7+R0ROf0fAH43jfxQlTXsmZtex7LfC2zx8dnSYdSJnB/dhCorAj/54avHRknA
8AWLTBwIU+PTYfB1Cu03VYFpv3WGjIbsNN2g6N/0JJgDka94HqKss2Pq2P7Q29B+
DIzZdYYCDJLZ5WBQf7sMDvLSRW36HbZqub8ipnlqX6XP8fADR/vLPqEotlJ7jmzy
AyoTi2vf+Pwir+l8mho5Kja9vcQ/YYJaj2qzdxUq0aixFKHhisI0EI+8bGlkglkE
SPC/q79/aQpp3vCtElE/tJSxe4jd+OlvZurcnD/XInlb763rnuqHS7aRs7hDLQ3z
JDXlbIcz8vnQKC4sQjh7d/caVQ9lfKz8CgQBtlhy33iaTe+XqGhwP30BfUbvMnPl
L+8PrCzE4kPReQdioR8zwQY43jie2N8E4OrpNOMMAmb5RDtOYhtIH2Wd0GJRxMBW
c/6Fqs+kx/HRoDWBbntX6750YuPgCfj9iXCNa2JVKHi0m/e4atiSfmUb+IdcavLv
eULVBlyV3Jm1mIysiNfTr9FKmY1c0p9p7GW+be4YAERMv40ZauIAyfzRdd+8X+MX
Ho7binuQXMDfywZuNSLzsO40ygOD+uARQAysw8FNXhXjYbM2COQDrKq70gjAYADg
cL0FLY5om2AHczvPdakPJ0yAKGkNgVpMCYFByuicspPi/SV7dOjkqJcvMlu02hby
zL+H8ET6r8a3eqX5XuWRHLfHXNY6Ai5zoIHPJWx32CwVn/wZxEdRjTXokwyinVsE
PswEjega1wZVkY8Aq9kv/LyePTeHJGXin9lP1KsFJJKQyGWYfpUTjPsHohzkiVgs
z5nsS0AuJJz6UlKIbjtn4SUM9SZCkBFAbUfwnSp56GJazm2iJ7zsN5pzvHHvGwCI
XJ5dnMgkIeXLnOPjrghKWBOB4aAshdLyRlcrm+9g6L7g8CyTS6vlSrS+mk/FyMOi
mKdPdZLrIMbGKraplXvXiZL4lFz6d0WZNxDEsuOFL700i5qavR0q2DMpZ1WpTX6I
b2REmInzazlzIXzHPE+r1cv5YJZj7Ge3Mbtqkazquo1f5CGnTwyCNxIs9wEMWCL3
meZ+rbAToFvpsiOD/PtrOxxjLxl+MTGy73zBi+Kd57pyPq23DvR7KhFI3WkReVhI
GSCX44LYkKi28vOBc/6KntQDtvS4VtAtbvNMuFCT8H+MekryQ7nbPMXEj5i4PJpx
3jNBW89s6TdNEjJlsaI8dF4PAJJNLA9Iy4CvmP7bFsnHRbbu1WAR86ktEOC8JWD3
I5YGLjGPuaoGx9IKQHeu2j3dd3QqvzC3OguKRcBo8rO5N8d60jlmU3/DNaMVdltM
tONoFmIB34xvj5Y8jHUF8X1sccd87d+beWEj/YhwonzycJleDwdmenE0sQqHck5R
gYCzDLoa3mGgPCwN5tRjCy8IkMet4CxMf4zjfpjVfijQWak0iz4nLLgS2oTR/HM/
0fnY5SiiVuw6GBcReIMIraYQsTWJzrqXMgcg/1MA6rB3sSzAgzyTQwLRrXvphY3i
0bxoVAckrionUCFw+B6L0BZapVUzS8+HQ/5bwYMAHwxNmtgbuef+udDDLKltYKwZ
UpyUG/ZqIC1BZovGaOlaSpXXYwsuj2VLCY+mflX1SdMPlB0hUN11qMk4mlXUtaE6
6JSUOg3BEpuMJnwaM2ttT1kuew5QlgKyPR0N2Udmi25oL//td7EpHcqiHD8jlR7r
AnjdVTzw9sCQDza8w6zdCo0ilOFBsHYSVV/pYAD5qBBRAN+KAWHEZ0w5RrPt7Fr2
3iSMnPAeevQfxvyVYCKlCUagAE31iK4gsuF5DHYl6sirXlFquRXGdhZOgMp/sahS
jX01jwLmK2+y5OhAvpkcCYfrfnnT9NaDFynVkpu/hBrMKOKJAQE4TezPg7yVDkK3
eeI9kpaBUVlYdlajXa+Jpe8tPI6x9LD3Cx2Of18d2CvHWu62WJ3hfu6wLQTOKHIn
0FCIDj5PDtgwe1J7i60/itvVLRMiu6cVobhGz9J4PbezT3ndEuetTFyWpTxXfbg/
w6VzQtCQrsyKuTy6HuxKOnt+RCr6XEySzYKAYTuoCjb9yajvH7DMuZSPkKs4kx3+
1nOpLTx6P9hMcXCiAyBRDYEOTOMCz0Du6LreE2Oi4U0eUSqMt1H9Nrak7BmxfKAt
Eln+WRqI/PTA39OS8gkNY7j7QFf9ClXTUDA26XDIB4ycS8+OkqSUr4ZMBWLE3xQv
WO6IBX97ML1GrZIQishBq8077vBwZthP9lYCriDj8Pxb/DPW1GQ27N8M5l3M8mLN
uhCKwUBrmvDgs4cWxhkc0BDDwYbW/iuXV3mKYPtJ3smFoo4HnesIFvBh3tQth2oU
G0llL5riwJmJ4OXHFdKQa7NzUCNi7+VOrcDiLV+7IvCkoSaax/VGxA6vlqH09G6U
WMN8/UI+pa50M+aow5zmvP1O5KNSA8Ov4Q7arxzsDsDV1zc9nN9KptH7VjOAx8Hs
QTVsKv5h4ciimMbXqqYYu7amUnd2stcb+fTXgM7QSS4HxkJQ74F3wi9tbQjMrH3D
qBwtXCwAwmojPoUDLAhiDYltn0+RzjCgWg7LIXztgGGdM/j3xTv6QzH8wiWqsefr
iIu498lkesTSDdEP+LqV6q4Wm3xJ7YSNk35uOUw1UGbUxLAnZ32iNhdzw54yR0AD
BZq1d6mmqpoJsORyHzsCGfNsFblWhU6lWi4+EzAUom67A1rT5SQvZrrbeZc7PQeP
Co+IQXLHr7ky3uolLDJHey+6zayoaWcfhaBNBWbc9kd2/Vhqf0wd7+ObXnZ1BWrY
4TmjaTEd05Md0QlH7V+nkN/gTDna+TiXswNyCaZEBupn6wMbuCn83u9hs5nlWmeh
CwctoU3uh4yuFgW6ri+6GpBnUy/fv/Rw1RIp0MwzxIQFN6tOO7EjLxAfb/zsvhTv
kBynbDhNjGWZ2zFOf0C2I0QRjeSai3MKdHJmiMuxF6LBiGK6xxCpMCKDVsAevHGn
G9Jus3ebrGyJJVRyKTTQ5danFEsppZbr3fOJ2qROkfZXtVh+SChQSJSsbWw2Oq/H
sVBHYh+4EVkc620QLDlEG7ksY//QIhaYd2mB1ZFWx+PT6PwBIdTIkraaSPYr9Qh4
QcFiUsLS9Pa7bAipLcXKo1xDwozlVYclXqbYgPX39hKt/UVdMCilWVUnfE6xyMd7
dc2/Wo1JCQli1oF+PE2v6HW1UPnw1dJe2eqPJ0ioul6c7GA7A8aYKYR8km39PNBP
0KO8ljqAXJy0ue3NM7Oxw1grHpvUlAVBfci9ZtXyojh1PnY4cmkKWvK8XaiOliJd
fvG0d7CxE5sOxu7p8n6LiD56zOTU2ZkdE9u6GwwABwFLrJKJlBOvh4urrHG75kpZ
zRWCrHka1jAgkyc3zrnwNeH7fz9R0gxwtiaLSupNw/Ny1KeR/xPZ4RBWHOFWNyl/
2OZEM2uARRD47/q1gIrXYsZ3wI15/kKzPLE7My+DCCFfnqqD0c6Ay5u3gn+dBG3q
XSxF2Ih+AeHZwVGNtr+hxDkaFVJ2iawBRM24zQauAbAs+iwZ789nnXWAniRBD2/0
gFuqw/0JqBz6+OkPKehzNzfaiBHVj1Rjvvulu4b4VofXGpj73yRGwxRSJFbPbMJO
oMze1FXEeqzAuxytxS9Zk4OQxUPGNFrH+IDylswQSZk5Z0KSLo26tB/VQGHSfNqu
6H1mFuD6gRZqiEOjr3HgJ4BHpi6bwRKFyI/DxznIyTS1DqWjOTY9ih0gz6Bo7uPu
DNSVs7vDG3W6xEGJNx0BlrPQJ91nB2/zHIAOpIHmCJ5+yuGy+RZwBx8UIf/aEAMs
avsfdZE3HC7S+mkpsTtdryUylS/prD5tIyEMaQO2uQc7X/YkWl1Q/gK/V85vNCls
T9GmARNsnB8YTHqwQZCjZS9ZzhGQAQSoFGS1fL2lw4f64FdTRdM4stRyX1srErLP
IaQVSMN14QAXFUIa2b21MVMv06AvBBWQ6dd0JZgtRwq3hc8XQjsgqnfYJ3rTjjZR
marNor+xWTdImcYqI0pCF6jPQMlY7Dk5pkbaD8h4EG+KcNFSbhrXNGnwB/0VrKI2
UAoLdycSy7yk4ChauCdWxQ==
`pragma protect end_protected
