��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�GN�Џ	�U��o�+|��������&l�Z+CY�G�u��\������j:R1hI���R�(upj�ɑ����߉bhZO���ƪt?���=&�zTü92�M�7%�~JU���r�W�לUd�$j���^X7��k%/'����Ҹ�{�`iw��Γ*��D��B�(��C��5���2��d��%~�	��y?��sz�ż��x�3V/G��.�z�?|�$�%�}�)��pw��E2�g�y�v���Z0�9�B�L��(H�t�4���$��t\����a/͜���� 
Z7T��s�K����Ћd�C��m�����{������ZOc�?�r��
%���0��,7�
@}k��;;�!gx`ͼ�8{� ��o����=�f!~h��k��/�,02�څ��{��Y`>ۡO�3^�PH����c��� ���q�+2[3�t�&̹C#f/����4/�p�nD�+���BX�Z�}`�����gS<�G��g���rц~�h��T������`�K�j.N�ܣ��:��ܔ���|!!��2^U�p4�+�i���Qw�oP"�y����D� ��r1�8�" {�����W�׽�L��u��:�˽-�����h�򫛉 �&Mz�s�{�G6A�/�����M��8��l��f�����n&q��B��L$�Z��p��ҲNN��d�}V�������8O⽂$gF��:�$��}�M���T�pc��"��,�(I������4���c�d�Dݝ�o�r&��q�.�(��'{Fi�wl���u��i�k����mZ�;5�Mԫm�?U��)�2� �5Q���)m#�
d�/��	 iJn���>��GG�*���"�ȏ=Do�ƶP^����{Cy�d����:�!l^(�bl�7�GCO�f�ԫ��t)ϖ4fV+4)E�MEA�)�P.�ګ7��Y�V�w�+����q�B�@ؠ�Ms�A�75ǯT�tՙR��Ϧ�$pE��"��Tr��đ��Y���LsRP}B^��~8��;e8 �26Wi�:���&�I�@�\�C�`<�?V420�B$��j��>ǈ��F핀n?_Pnh�xɔ�(.��&�|���L�)��ٗ���Zo�k}>��u�	=�l�k�"���:���{L��Qr8��TCrv?>#�޿�.R����W�������5��ҫ��(�A��5����I����-\ʹ��dg�:���9"��!�i8?�O���:-Ӡ������֋p�pZ�͖�*;w<�X��x�7�L�7z*"��G�isI���}Y)K��eE�����x���^�t����9Ȋ*:��X�D'�(y1k4�'ͻp����,<�kJ�-�k$�}p��$'�+3��şh>�� A�x��n�$@xG<��'�`�,v;M�̝��̝���_���$�~��TU3O��aYl�NZ`y�'���`�R��ϒ�I� �ѝY�:�����_��4��W�c��E�AF���]�D�� q�(>���D��h�� ���zز�R}��@|'R��q�\��^~E��T�l�^��<;����W6����Ʉ����l}+���k�odnQ�'��C#3og��/M�ʪ����*�b�	�T_���Ȍ:CSR��y��g r���*2Li,px��m���ػ]u�_&N�SA�"1��r�0��?*�N�6�mH`H��?���+>��#p�zf��<���*x(��g�q=��>��� 1/�oF���3�G^�]�f�Y)����[����,�!Y��\��6a�S.�}Yp����٨��H���;��2긠�	�RC·
��������
��P_�E��$#A���F�]��؂���D��No��[{TY�簷�DF��i�iѿFq��x�qr�ddi��lR%&��#�#�/ʩU�y	��x�!]��j��(#uի'�C�\����L<���ڰk�Hڿ�j!�*T����<��Lv}��b�p]yb�IE�g�ָ�v�K� �f�d��!�;�7 M4�߉#�t�_�=��O��7 њ��
Ru�Y�;[��=� ��=K���{�A��ͳ��)z1�|aD� 1�!ոa��f�d���N�(;h %&Y�`��{���xHM��g^FUɴd�Ѩw�u&��8�{�k ��,��d=y���u�ޮ�u�̀sH� }�*Cq�$\��g��rIߐ�h@�|9֑�/�=���kNY�>���5:;�P@s!�x���_q�8�Ȧ��uFHpQoHȱy=�:���S&�k]w�ˤPA�a��_�x7x�wJؗ��i�������L�鐶c���^U��UmX���~�i������SR��71|���^z�y8�Z魈�����^�ME�̾��A1����\�s�9������������X��I�נ3m0%���
�O ���͛X�V�`IC��Ǒ��j���X�L.y��g@n�:���I��@2.��
C���K�B�ɍ��Z-Q�4�(-��x����3�k���B���@n,��f(�0�$8���̄�>�6%,�*b�
�P��ğ����ֈ᜝<�ac��:�h�e�(���+n�o��s����gZ  jS�
5�ë����c�[)i�	�^�? x��&�,��ҁA�,��l1��z�;����v�%�9�e4��'`�̂����wK� ���M;���U�JM.B�aJ
/Ak�Ȧ\L�sXa �'��o����Bbs���kn΍?фI@�u�J��R�Hw8�V%[H���8�皕��m	F������f+�	Z�'ޡM0��F���4#�1Iq�b�>�Lq�6!�ގ0�Ï��uu�fx���m��(H�	�K;.4a��r�YP��v�@�����Fa���w���t�C�lm���"=�&��	����(2�<�Pgw;�5 ms��?�9Y������/F��H�m�4g�=p�%�$Jr����_?G��0��z��ݓ_-���v�\TY$2�� ��U KFN�}!�1��P�'����k	��>ԗ9K�@,���sa�N�"*a� �*��eQN�ͧ�(� �T�n
ܺ��(�?����מ�|�o��В�X�UR/;�*���*y�B�Sx�~�o���~��"���WeqDW}�*H)VF�@k9�𫇅���Ū�8췽S���m�O�q�����,sGo�&��mK�9?T�6(R���F2�P�o��3�(toĸ �3������0B���B󓙍�^�m�`J��h8ˇYq�H�1i�����G�~���]M�C,��'֓�dXs"XA�ؽ&U�ң�@�5`�'\9+EX�q�P"�D8G?��7��ͼ���u�4�3�{?(,T7F�}X����ϻ�Յ�֢N��5��y�G���[F��Xm�|$�����n�J�����
�ށNtI����n
>����:�^�u��+��͐�}$�cM��V\n�����x�9���qǵ��B1��&x����t��[�'>����|(�p��w@=����;�-#O�,��z�%����������T�oE?�k��f���]4ڪ?�o��pjDc(��'D&2\�2�]���
����x�<ۧ��#���Bs#��{st]�E����>=���f�L����V/"�Db�H@{��x9�d�y������0 �1W��i�@��޺ϖa�E:�%ګ:���3D�1�ތ,�т����Ae�,K��|s�/d�p�VR�iB��Hd0�v�l����@_~�~���f揌�����bT�(p�.V�����a3��#���uJ��Ǘ��*��
A�H��.��O�{=�o#�����q
�
x�489�<�v��P�ز9?n��p���i��椕�OBb�L���Bb��{��t���L�o���(o���170{ގƳ���N���<�	O0od�}Dr�A:�F�/���w����թeD,�#��*P�+F=�s/Ԭ�����������pj��T��Ʋ�U� �3r��g�d@�*r[4 OB�Q�����e����?+"6����+5Ho)r��&��?kLF��)�8��c�X����Nw�1���t���[;4A��f*	�N	l���k�4o�B�;�M�7I3�y��rg�T�\��
����Y&�a�J�r�0��?ٸ��2��`��\�Cn����[O�LKMMO3�I�J��e�*�\J�2��څm�5����H�"C�����aqnU&A�����򟷡�V���N����'@%��;��̙V'q�n�e08V$�`�m�-����ґpF��.G���]��'���:��S��5hϮ&�F`��wsޜE��aT�H!d��ĮۓJwH4uj��֐��R�\J;l�����؆�B,X�d�ݏ������ꓚ�Z�ͫ��y/6*W�-��iSz��\0m41�o�}OD�,�? 2�8E�I/��a�Yőt)�:`>��D�jb�xj��C�x��<b��+��6���
�N��rwb�)�S�D��#J�9T�+�ׯ�E�������}��Y�Ncz�� �'x^zثm`����J���VP��/��&�bm�_��#�B�Ni '���}F�e*l�\J��+(�{$.Va� �H���Itg�:	��u8UkZEp�}�>�U� �Do�e��R�P4�r� i�q�+��4c���r?/d����8R�2���~�I��y��#4��`��+?@'��d�Y���=,�i�{�J¬��� W��F2���f7��8�#�e�l�O@
7V)r��=f��ʅvM���o���gZï �b���TF\����I�>��wj�{ЬS�[��)a�}��T	�ׂP.��{_2�����%BKM!�gD%C���ǋz}(�v�t�>zo�"�`��tˇ��)N	�T����ϓֶ�t�L�#��"$�Z�K[���8���$X�W4���/3Ja��j�/Bp�6�-��!?�>��@��'���t.�A>��Kb׿���M��O��&�ytX�W585��g�\՟���d�t!՚c��bB:{�ة(w��|`��N?�55�L�+�����.��1SN���gV�>r����G�1��R:{��쩮��>�uDe�;�+�_}��	�+�M1����1���05>;sϪ�F8���e���'oV�(�U�Q�k�xTf�����p=}=d�Z��Ug�v',���b�������L�j;gQ;;�R?qY]/�h��B���S��:�� ��×P�F0ALq�b�F+$m6�Kr�۶ݟ6��8̮Dڣk����L6�:1�P���oY���'3��u	v�~䂃��n�3��a�-��VZ2zʠ��#o<�x�C������u�
J�$"F��k��L��=��T&
(������ӌ�5f���cl����`s�%�� ��u���]c
a�7��GJ"�hd�ie��/.'?�Q2��5�zo�@M�����W�%¿sX�OW���Z�ߏ�>S� ���@O����<�a��M�B�R�%�Ejja��Pjt~��-X�Y����!4��g_�Ө�~|�N�
������1��'Z&X�=$J�Ќ�h��-1m`~-:4���85�������}�#o��H���-��ޙ/��ں�5�L�(�X�n�l�4#[�ճ��()Mf�:[��T��:`3wx�������bj/���>qu�
;�9q��Ǐ������Z��c]��B���M��Ί���oT�x��5.\���'�Y�|�C@6�����ѰIU]s4űa��$kU��ܪ����^c��Y)%LU�[�@,�ߘ���t���d]�o��n�����VJ�Ur�b(��S��[K�M��[7JE(�*`%X�h�\�@���f���-��&�_���g�-��}w��:z��?@��N�p����3������9q��L�D�f�8K�����csk��TE?t��[��;��1Y��k[���z�m.B�ڡ�8�����ޥu��=�Q���������b�b����VO��fr�j��������ʅ��r�h�V,��zOq�=*w0����;�N@����ړ��.���ӗ/�_��#��]E"A^�)�Z+���K�^Ƽ��F�j����°������ �,��Ki{�duv��{]��&����h0�Oז��|���I�n��V�ϯ�����u��_w�ҌmjGMdY]';�H�Gv��b��V�R3e�@wh����I�6�.>��~$������HnN�w`�iiFH^�S���A^}̈́
 UD�k��J���R��GF���+�g���T��?�8	��e9n�-/���7cd�K�B��8���rQh܂M�r��{����vMT��/1B�ҭ�/���v����Q�Q�%b����l���V�;Tl������>yb	�«1`se�|�RI}�U���7�r͢?��Z�妙r-?�d�+�F?Н����laAb�*�X�)'��-Ҍ�i����:�#m�[\��*Z'W��V`�7\u�_�v���:[E��.��q�{mP��"�����X�g��������/�H�pW�yl>H������W������\�������ӭԙ�@t������r����gMbH� k�2#��D<d���K������ꈯ1�̥�UT�_a����7��#�T��5���l��k!��z*���3lk���⮩�W�c\�����JB��u~�Ү����w�Cl3��cf�D#�"c��Q�M!v���=c�\�U9lp����%�XL�k� rm�����eT�;���Whma��`u��|���LU�˲� 	���3\ /LMDH��r��Ƀp=�D�g���w1��ʹ�ח4�ӯ����)���ľSXԠiy����F&����d=�\/}v^���9��;BS��R㉠2�pX읓�M�䅫plF*2��	���b�&��Do��h���h���UXZ�]���t�yE��Ň&ї�0q�&��ƃN�%�r�K2mul��$��%|�Z�3^��h�y0G=�i�#��w�f���7A?��),�X��` =dG�I�5eil��}���� A�4C��OE��:~���=5R{]�����׭Mҗ^3$7��[�8����H:lf�q�N���k�Ȗ��@J4~�����"�1Ï��.�����9��"�P#�į�;��TTܠ�ĵ��i��ט��թ�LI|,�b>�8w\���f�v�g�������ض�C�H7�&�'�w������N,*�=kp�~RI�f\5ุD��������kį+��ˏ���=� w;]0��<A
��|T��H��$rSɢ�r������U�M$�� ��F";{�	�'�ۼ���1���_�{y&�VP�j�N�A��U�L*e�U���c��S�Eh7UvAj��{&�玲���D�����®d���hG䔺E9�b���$ʌ���C*}�Ƅ����,/�	Xr؍P���}g5�ߝ/aI)�jx�W�-�=�"��Fr�����`IJ��5�tY ʹ���V�ũ�6��1�K͑ �V��̏F�P��-���o�G����nv���_⡌6'���W.0fyG(]0ߓ�g��O-nҥ̰����N�F�ܗ��T�mNख़S`�������L�RD��2Um��Q���-��|�lp�kTfİJ����By�Hzۘ~
էS<�6{�%�<�$Έ0C��ϱ����C����1��A��Թ�����6F)�@9Ē1�v̐���/*��z>o�����m��Lw� ���,��5WYpKC������b�a������?�`$�xs $z+q�NX�o)�IG7S�:�x���}�I��f)ѷǎ�tocPl�4�)Zѹ�jt�H%N�K�KM��x{���G'�5��h����jwv��Z��
{a0��Y��%��Z�ՇM��[�Ҥ�ƒ$y�d������+��H_9]i�<3�?��f���2c&&\(ϰ0�� ����	]j��s�^#���4[�&������]�m�%_�(E�-Ӿ˥|�ӹ�#��c���#.��iZ	ʍylͶ�k	��hRZ��h��
������1�B��k%�;E�R������ž��[Q��Y��ݡr���Y��y�@��A��G�:3�W�NX���k3�O/��8t�9���k�ဒd�a�N��\bEH�^\CV�Vh6#irD�� eE��xW6,1 /�N�_~2f�>��F�S�8/t/�E��T��+�ߡV���"3���RN{ �lI�����*Ӡ��~���9�SD�V�{-K����St�/�%�$�.�G����:�w�L�
���-n�j�V��opcz�'��L�~�y�ǹ���{��5����L�Ȁ�����^iJ�R�� �T���$�#��Y���R9lD�ĦQd�6��n�Q�����@[a�?E|��hιJ�a#.�q���D&��nZ�P��Q+A�#�=d �~����X�ן��B���|ʬ�6׫n>��^�j]=ܝAm�M������-�o�+\�ovB����4:Ė���
�Ű��T8��g8���:54�n�~A��r:�E�z�]<�H�v�����z�Ҝ���f*��]%U��@�<��&���/R��h��Ф��K���<�۞Ǚ��*������-�9~�������������ElA0�H��5y~��-$��#r��Cd�%ةT�Ev�H� �/�$��?�<�,W� qݲG�-Q9�ҥ�4u̱I�v�J�R��wKˋ�nx���Bb��"v^���I�J��	I�(�PC^-j ��}N-��(G[���
Z��a�2
"��8�ȲAd�2}�+��e�
�����G*V�I}":+#6yD�p�PT�U#�۵LP�ѐ������8
N���k�(=o$�oV,N0���C؇�n G	�a7MXrd��"-��0=�t9����&����W�x>�W���ۆ��"Ltf�I��U�,m6�U��n
�l�����g+��da��j�K����	�������^�'�I#�p�!8	������
�uV��|!�����=�l���3!C�/�z�ԩ,`^%��k�#�	U�WlF6�m:d��xLy��%��-�������"6 ��c=X��ϯ[���ȇfJ؜��"m�=R�H�����#8�:��h��w�h
�����/ꞛ6�!�O.�98�7��`���e&3%J�%ܮ�:_�{:��C�Y�RHhf#i�p�T!�љ�F��g�5�)�Ōcg���-�U��5�L,�&̨�)3���)������w�I--s^�Ԍ�o��ΐ��?�ⷊv��kx��'�� �u6�B���(�h� �e~���u����i����S��ה2�E��!���Дn�:\�7����k�}��_�v�\��f�4*Vq=�YnQ���o�2�ܖ��\��ill4t}~KҼ�M
���>t���Z���6��l��p�Dk"��ϓM|(N��Ȼ� �@e���W{=�90 ��FY���8�)����Ι��q���9	�ϴq�WDKR��)	�Z-���7�\���^�����;��}�{X���m����1�A��\}�^�L��A*e]oN�7^e��K<�L�1�?�uZ��)A��T�(�����f�\�lb��'T���J?PXp����TQ`N4&b1^3������	vCQH\
�C&���'�U-��F%�?�Ipf��i�և��K��\���9�994A-���{Ov��e����m��(�~��ՙ6Pv���p����';��o�"?�=^0�<	�~�c�U�ޤ�	j�%��Ǹ{47O���j�pO��P��R%�'9ڲM��{6��B��U*A��2ta�y<��}�Z��������K�^�-U�Fx���{M�<�� sh4��.T68�l�GO��c��v�sL_#$��\�e���z��*�߃*3.�!����U��a��بU"?�t�q8�R7]�Q8Wʹ�mn��%�p`a`�M�'3]�v��V�ɱ��sy�S�����TtFDX��������5��Ֆ��tTyʗ[����"^�$3h:pA������-��,�~E��tЙ%����?D�D���R}RޯsWG���s��>�o�c���[�X��=��ݡuE^���h�fzW���P�c��0'�Xu��.� �7����b�R���y�����"X�0������Z"X�,��Ԯ�����&ё��ui+�0Lm�����;�,��I�J�5�Ò�
��3����7dN4A����!����S8�� �k��j�Km(-ҕ���B��ʋ0���XW���\Y��#������9T�i��#�[ۭ�aX
���;�Lt�C/)��7�鍜�������LmKg�Ҋ��JD{����Ӡ_̏M-�N�,v��\P[�P������j�Q���P;\���eb���K�<�$�Ry�Fu1�����Sb�6+��
-�b�l*�2������%� �]4������D]�ń�L���r·45	�,9���[$U�A\t�������p���;mj������Z��Rs C�Zr&�
������ 7�Ԓ�3ٰ�ϒ�Fn�Li ���Ļh�[�s�?���҆�ws$�-�{��2+�9��IT���c?���u��O�5�iE��]��i�~h�[s>/�x\�,�u�=W��;w�}��E���y���5@"�Ы���i�$�o��<��80/�I"L���������=nk,�Nn�
!�|�J�bk�S��4�	�+)��N���d�� 8������ԃ,�z6�K'�gߦbM�k�:#�E��~�$�ƙ�*>�6J�砇Q>��~��#>Q'�Ùg�)�*X��&��M ��m��A�	�meJ�ұt��(]	�����*8u���288:�:sUjP\Oa����O��8��[���2R�+E��S�?�w�V9�E�E���[2^_��P:���JH�t�=n�K�yW���k��GM�m��æ/�4�+W����Yeߦ��ѻ  W&"�^���|j6����osr�m]�U){�{0��+gf�,��S"P)�Ek`4!��>�E�w7T0F�2���J>B@E�wu}�^��7��-ړ�z��SL0X��D�P?K���,wb�%�2�c�wZ���"�B��G�H�@G�e��BDi�o��$k���.W|�<K�6~�A&sF�#�V?o���X�\��%u��΁�wR3� d���L�����h%������ܤ�(�~��g:�����&ý�������a�d�?1����pNZf���H�%�:��]���N����ܞ�S��0ق�i ���cB(=��,y�j�O_��nD��W��`�e��K6��H�����M)��Q�|���L>1*�[�tF�Jy����J]@y�p)�ޢ���"���Țl*���w�=)[�ޏf��H��%Y"pS×L"}ظ��KV����˫�`l�)�'ӡ�Z�>J:=�~LU����H��)#�m'̾p/V��%�<�SN�~q���[��¿>�x��I��Tz�����n��N� ��ΨY>L����?l���c>h��r$[o���DK��Լ�Y��eݹ�pƃ���,I�Z&�o����p�ƛM07dU\,�M3>Z�� dE]A�x���FO%�Ј�8T�1�����OhPlޢ�p��1�{��к�NW%����
�\���Qa��)#�_�@m�t1$�ØP���_��3��[��1l�5^��Y��<qP�0~,�]4���P.���N��;�U}_�3�9�5st���g����2ݝ]��6Y&�f��|�ӕ�
����>	tD�܈�����Z��S��V�>�t�Rٳ����ϰ5�F2��f\�L2����]��(�a����zq�i@%�^��Ǚ'фW������a)��v��ax�Ѿ%�����x��;�n��|L���(M<cM~�ꈩ>/��,Q�%V�Ѝb%�)�L[ >�
a���*&ɗ�ݲ�ppq�o���L׭�)�q�U�E1~�v<�؍�_)����	Q������Irq���#�I��@�L ��G�2Ǔ:JjNw���4����b����p�y �S�9Ih'�W`�xc۲��j�>�eGR�#(��i��ŃH� `����b?��׳�$*��S�c�;4��7f���7��;ٚ�����WCl{�ڡ���.2������iE�u|S�GW\}������SEy�A4T`���pn=�r�Oh��X�Y m������%n�{:
	�1@�M۳�j��?짦��g�f�mc����-IK�BC5�n/+Ԇ򸴄%u���|&�6#�����򵶄������4+<�*8�	�]���`$�D{&=z��^
w���͹h���c-��PH'�k�w��&OQka��J;�.
�5R�e<@�ؠ�)#�� ����]yy��@KV8]����#������>Dg�;�;��YŔ���aLf��{Ȃ��/QpǼ��
A`N� ��*���9��a&�4΁@�	Uv�	c�͈[�m?�&�h1��Jb
z��MJ;N�_����R�HJ��6�!��4�_d��Z���+�~�&��r:��D䙦�K*;�˖���$��f$!��^��R�7gخl�f�@���B���]F�k�&�q��WM�$�㈟�6�
~z!� i�ǯ�BU�R�<뉵�l��_�ċ}5�^���b.ԿKA���&��,�1����݅}��<p����|�S��-.�ҷh��z�M�����|�j�`7-��|@5��HP���/M�ѱA���O߯�
8��Ǒd�ZPm,D��',tV�MEj����@���
)*�~�&]� ��H�h����bc�͌��zj*_˨�Q�oܒ���Ӟ5 �]E��?�B̶��X����wժ�>��A˹�֎Zmc�>�>�ʨ��o$�`����#��^�����p���}�̆��U�l�<�*�yT� ��v3yLB��`c�z��K��g}Eg.�B���xsx�h~��l9<d<�Y�j��5��.&�u���@�L(��)Y�ho�6ѻ@�Ϧ��Ʊ�o��*`�S����:(�'+]'= ז�u� U��6(���z�(��<%l��Qe���!������+4_�r%1�{e��H���I׶�!)v}��}�Di8��zs��U���v�p0ޯk��Ɍ���Ĭ�h�\� �0�>v����m���e#K.R;\+-�	�X�X�3���.<ՉTE>Z����L��-��h ��.��`����'h&�s�ɵ���D*�=���р���q�4�Ndm�1���.m��n����p� qwF^���
}�R��4�.w�"O����n>4ak��l^hڑ�[|%� �!�߯���Meo�u�Q��G� �����UI=K�
-�v+���k��M1��%x<I��e��ܠe]���kzT��'s�,�/�)`�*�n].RZw�IO��M}�q���c�0@1̴4����?raafx�t���z�v�vOٚXz�Ȑ���'�.���ѣ��Ý�T�b���'��!�o�d-���0��dN����%�%}c�A\	�PJ�Ts8��m�t�^F��g���ݍ �ͦ��a�20*��"{�����R���Qov����q �R�e�Í���{;ɡ�ij6�UN�5��v�߲࿳
2r��A��� #۬~�@>��f9�Y�Rӗ&:�+m�&/���`��\6�,��؏��!��< �zA��xxw~U�<^9u�A �h���hjW�N�~~[�,{�=�R��Fu4;@t�zv�(,X�ԍ	 �3�
�J���7>6�1|�w�ͬ���:-����%������,��V���x@��Y�KLZ��C�{��!�^Ok��	���Uq!�Fv�uL��O%�L��ꃅ���dR"��߶�O+��FҕH��`�M�c�y��ѡ�sX"���$}{}>s�
�q�|�����CA�9�e�T�d���,./~容ߺs�f�;�<�y������qq"o�~�9x�n`�kHV�!�&�����z��8��`r#B�oP[�D�ҍ�с�s�^�����eI�T��e���I�FO��~���|Z�%���!�x�y�/�N���5N-}��yp�/�!&�<�5��7�u�)�n�r�/C#,�k� ��}Γ����>< {�	h�˒����<CA�ȏ��ۻ��6$�pA_�QY�R��]�S{K�Z#��h ']S�_��ت܈��LO���0�>�����ѳ�l5�ê��ƫ?��Il���7�C���XA�w:w�!�T���LS޻+*�ƞl�A�t�d� 5X(olC!a���o���*Y�J��n
W����}��L�|oc�̸3��!D]��>�*c�z��U$�R�n����rL��۞�K�E���KR�:)�IK�L��u�d�٪�Bv��k2���!��!b�Jg��G�SV�����D�-�j�8 �N�նZ����{�Ȁ
���6gb��y�C����f��i��+�N��-.�+�/�^��L\*I�'�a0�z vAHFf�1*\��b(g�}'~pg��p�Lagmw�]Y��tR�.U�,��=�%�	)l� J��ƽ���ߡs�6���v-<+���o�b'���W��V#h�ҁ�F7.�����O��|��@�~��c88�b
M��=�4���}�g�	U��w�뿝f������P�J)��]�cقA��
�2�*�U�Y�y�>�0���LW;����%w�5
({��w����{��4��c�St����̳����KW�s0F$�Wӭ��o�d�<���ܠ��ģ>�e�����na��Mj#��a��Tv8K,g�9�U��]P�l�-
?^�)1�.Q<�^���l�"�}�tR�Դ���^���|�?>/y��v���� Ii��v��q �h�L�������D>���R-��{3�NL
�8!C���~��o���§�\�KA�뀰��񜩰u��"2!�;��1�2��&ӷ�cl�vu�?��l��p� �o��VnƂ8�RB�j�t>V����v{Q���0�� �C[E+������k��5�a�Z�M⋏��N>�;��6��^^d�?>�����%(�nT���'�F�����8ω�s<���)��,����S$��wh.�Å�ȈUH+^ѱ����H��x�����R9|V(|"#��ڧf�H��@[�3�;�kK8�GOv˴�Q83dʀ��-2d�丒;�G�^V��~�f�����Aw �n��A*�|�	���ʉ�7k}����pϧX潟�D�2�E�7�J3e�����m=�m	x����n=�[_`�ݳ�FZ�f�
�T�A&m��Vd�� ɐS����}r�߾� 3	��4������;IPL>�@j[�O�9�Ic�7�������	M��L����K��u�1�u˞��d|q��)f3����>A�R��hv!�*�ig�YTH�R��� ��P�)�TS��Y�t�(�ӧ��u���0%��0ꚾ]��	�6k�z��1Y�ͬ�l����3t��#&-�d��l}�UM��)x$���'��{$�>g/a���aٟ�ߴ��8���?�����֟!nDd��䶌0�}�I��}�N�e�����Bw]K���n9��tOr�haa&���1��z}���q�ˮ�c�dW��P�D� ��Q�P���^�̡�C*_lk�Sqwρ��{��Ͻ���:�]��o&/�O���c���EK�zZ��t�_%���>��lf��o&j=����_�a�o����G4���j~��9�����YOA7�w�Cv�7Uk�EC�K���$��|<��oǦ����Cf�7��1���Z� ��_��C�|L4?����M�;i���p���D�2�]1b�TO�.�^t��$�noCi;ɬkf�Hs���S�)o谨V�6᪎�m_��>iN�%բ��ZX���>j�Ȁ�K��AIY�����n��
��ll:����!������}��q���ȋTs�8�,O�f�� ec*'����s�G��a�;��q=S�Ȧ��-��įg�Aǽ���r�+�U0m��N ��8˛�'H��d�v b��B`�`��G5����SW�Zb&'#�_ֿ�YE��r��B���J���m��ޒ.k�i�:F�JbϠ#BІR�\������h��"��H����O힞����ۏ<<��QZ�æ��EVs�[j_F������#�E��^gW^��/��ʱ8T�@e�Qχ����vEqE�袘-�BNS�U��T��z�4C.���l��(��Z�� r�g�[�U��|����	X��X�\j��]~��v�~�Q�R���n@��-�
58=�6+�ԝ�i��2h�3������t�o/Q�	��h�C�_|�}��2�%�p��t���zR$0Z*w�?�ŧ�˼5��8��Mm_�?���So@O��~+�m!<���|=��$�	���7�<Zg�Iȿ�8U�$V�H��֋,���Pq���?ح��խ�'M_Z<���(i ��N�&�am �g�_ݬ�yR�3�����.9�gp0�ݩ��#}�f�+( &�@o����������K��ü��`EG����"+GR��Ì��$<�s�V�=:����W�_&
$��I���V���.��u L���El{H�e,����)B���4�<����w8���Xb���.��S�+)Fx	Q�W)F���v�%��X��C ������w�Gr Z�Z��ie�3 �G�V���E͌�Gt�|B���頸J��{���u�f^���:�Y'J8J�~� kL��Nh��K�j��8Z�c�=����1��=p�az��wInҔuz���_���R`
�&���LJ��U���ﳄ�� �qtշ��b�g����; )����m�k��.�� ��\cڊp�L�Ⲓ�߽��8"D��R\����@3�FlĆ��yk+�S\�w+����ዡ�M`��x:U��g��cT�H,�
xD,j?��s�([Q�0z��J��q���A�Ϟ��,��������[���*�VA #tA����Y�j�ebݾ!m�{�"�n�cr��d����r���t�h��<�>
�.���Gz-`A�0�XOrٞ*-��OA��d�n��x��{���⦟�_�y�{�^7�߿'m�w�ͺps��m_iKUWg�1KYo�q/��e�<YuSm�XK�`�i�/������g��m���zVl79�G����v�m�캵Fո����Y������4�})��-��a��-4����D��A��:����{�oDa![���ą�7�����w��a��N'�|�I�1}tE�O�� 8�uϺKVe���?|�*��KE|��Z�%��J�4 �:���u��U��1	{f� �v���z$1+S�w��Ȃ�J�B�L��$��/��:@0��2<l)��E��ۏ}�RT�D���}���]�)�(�Nno2�覣z���[
��V���g :�ׇ�[�,���[=�R^����)�rk������oUd����Ea�^�ē�r����1e|Y�^���L;+�T���JF�ciT3�s��x�a.s�����L�p�$�ք�[��ʷ�p*F��!�.�f_ʛ��u���"�Y�+I�J]>���pFީ])���*�4��{�bA�-�� _�|�b�4��ILi�A[�V�U�zQ�����H�r8�I�;a�j�AZ5�/�kw���E$Q��fL�rᲅp6w)��Ȩ��K-a�{�H_8�� ��ӋE(_���a��y�c�����{ �ψ6�C�
5��R=|M�6�7
=f4䷈�9�s<.�.�n!�P��l��Hk�$��K��t�Uԗ+>6�U�k H�)�u#�L�)�U�}�i5z�/��0�A�C�k�(]��1"��j�P�ncOh�̞n��eW�Qì`uq��eل��7���6�nc%�z[Oǟ�{��U}OEʫ��Sz��,bҊD���0ߘ�~����Q�mj+���fCe�R�����HbY�uם'�;�I���(*aj�n���0)oJ��>вN{:��@wbW�6"vUY��m]��x�#Y#/|����E��S\�|�_�
h�w��qݪ��y7Z{P�&��1lȩ2]�23��{氧s*��pK� :��FY��a&v�V{n"���wP���
��u�V�������;�����p�ʅ�H�����s}sf��ZA��?�(b��I���C�=C���z<������H��Ʀ;]�&�#�@֊H�)LE�%��o߽}���+M����q�F^rF���Y|���.�,�0��J�^c�7�%��|UA����O�N�j�1����y�Zn5m����e}"���;�/��Z��+s��U�(��0������w��dw!�Q#��CV����ax��,m���
Xa��#����;�JQ�����v������8�ҩ��& �����ї/hN$��%�B��"-�#�2�M=wγ�4��ף�F���:y�����&OV�h��9��{�J����ɰ�C�Ƙ�?_�=�c�2��(~��r_J��p���k���=���jp��@�z��ޔ�؈P����H)�_	��Ż��L-^�Z��:��Q��a��:�*T���|Z�˷��m��P5L��:�� �Sw��(����8��hU=~��� ?.� N�Rzmb��0Ǳ�%v��3��>,�,�����\��`-6���g���c��o�WJ��7�E��opU��=��%��ү�­*e��?kE/���*��STj�|ۥ+�6(>�7��?9��tL�c|��G�������=D��^�m|�q(4ȧ���x���ڊ�H��1�^['ciRA"ւ��ڻV�iI��K4���T��Yij�NG��~p���#�d�SRJ�d�q��<��V���m�h�d	����>�+>8�����|�)��� F�գ"s���v�h �4s�j�ԋ��C«�g�Z����1��2�[yvV	�׬��b��)����j�}#v��ۓ���6|ܨY���E�Q�!$��C9L��^���p�e�����HK��r�R��~�"��_��A]�%��q;1J/��-E#�L3�=���C��H��)����(Bj��к��]���]�i�.A��]=L�p��QZHP��/ь1���Sj����A�fC���f��Z�&�Ɩ���$�[�<�+���~8A�9�lBUrv���@�a`�D?��f&5����������W������*1�̹r&��g�1_�d/��}�۞��<�
�-�򮹲��0��"�%G��I�Ǣ��<[hN)ت5X���E�:�{�Z���6Q�՗�W�&#阔�f�y�`���o�=��+����A���`�=
=�pX=�ֺF^��0S�p�קb�铇a_z���Gŵ^��d�9�p�d��S���tK�^����g��"J��r�e�Ą��*��.E�Q�����Q�m��Lk-�����Q"ͮ ���3&��L�a�M4��y��P��]-�A��lմ��|b�i��Z��K3g��v�7Y���Iwt=Tnl�2$I�t_�tÈ��NX�A[����NE��s�_���_`��{/��a�b�jF^���/�O�M"<׵=�8ߓx�h	�~���k��`���U����;��R��&�_X'�0���8㾃A��6e����W�9';�C��$0<��������E2Cxl��	A�^j��苙L�v�W��y�ELs<��I�dM��fJS2�bk���|�=y�h?�fsO�Ä�9��k0�<�ok�v�7淂~� ���_��Vܸ���������pn{teu���M����� ���6�&pʒk8�U�jE�6)�c��3Ą,��<a��Sz]�Ȱ.3���g���M�M<Bb��g�j˙��DV$��-Lܺlrz���a)��j ���AhW��ʫ��I�ۗc>��v��u�M���|�0�X���`x���5P5ems糹����v��0�[���ʲZ.���̕�{̀"9f���x>P!�e��ZI�G�b�+�?:u[8R�o�6=^#��U�yL͚��9U��K?���y����{���$��i�l�Q%(��Ã{���!�hI���6��h��_XB<ሦz�3JTs��E��B���E�2�Ǉ�Ra�Ɂ�ܒ�3q p6�kT�;��?CuH��}u$b�b#��ά��� �1�����`�@�qD��˜_�n�;�����J�W41�^�4^�e1���w�n���]�Xv����q�u�A���D�#7'D�j}SBE���]Y�D��W�愷-���&k@!&�N-v�u)���o����9�~|E���bZ�_-Aw\K.f�w�%ʵy��8��V�Ř��6(�M�@T?�c�\o�%[�ZȐí\���rH�8��>g�|�֩S����=9���k��n��� !\��e� �o�R��X�GHݶ��&�C����{Yޡ@���KY��=��귰�=q�5���m��;�3��7��X��X�}��H.)�Qi��>"Z�w�e��_�\�Y����Ǧsu�,�qk�pR��󮈄'���szxA�����NV8�\�@�k�� �b��˗�&�>�lF���D��[[Ъ!���4Ieǘ�k	�&J����ә�|��n���31!r�4�,������9n��i�&米�J�^���,��6T�!u֎��C �(=���h�M��GG%��$�D�	C����F]�%�n5��>�eNa gl���+K�<S��lsѾ'������}��9��q�!|_���^;�Yߞ�f�)=��a�q�`~�Z�a ��\��n�m)��h��Y�	d����dÑ�Wq.K N�c�U�q��\���Ms�Tؿ?���Ϊ��J8�u^���x��fzX�P�2�-ȋ������D0���S��G� p���Iݳ0�\߆v��LK��k�'ݙ������jnX�?�)�A��f�& U��f		�1�=��Jz�IP�`B�rR@�|L�h����̟'_�ɗ��䀣�I��%�Kq�ym�� ~��s��u=�n�G>�fh�^�?V�(PJ�2���K����q��4.y�i��u����)X�!���d�4��S��ϴ�-r�-S	
�b&���o��;����0S�^���s�?>���潽�L�-�\�f��;w�p����>p���_̊D��*����yMll=��6�1t��w��qeN��{�������p�`���&iY/���>�ol�4IC�lue�Q�~AP��mI�s�2`��W�u*�o��H�C�j+�a@�b��h���g���Z�b�'�ݻ�t�z�y�4m�P褛��^��h՚ ��l��%��5f|�s󲏘Lo�ԏ)O'����>83�����0��%�����f��Ϋ����K^�����r���8�����,����������<���}�W���5�Ō������p�zP�z0.��4�M��4��^�����M����zS]`g,kM��o9'h8�`$�͏ j̙)�1��,:DXǭ$X�c��"{sxNri�Lv�8Y�щ���ů��p���Th�����-��oa�z�E0��p����TY��B}��F��ʽM{<LT�FS���D���D�گ�J�X%2	��Lb�w���*��ٽO9�����Q���i^�`~Y���-�K!E�(hJ�襀�����i�8g����Z��r�`���`�>?�Еy(��] ����F��k0�E��iN���p��ݞ�h5���:r a{w`����RY�/�������1J��\��sg������E���&��l�R�0}(���q!N�Tn��S|�ɧ�#y����~�lIͿ�MVvr@*�_ߒb�ʋk�rz[��,y�����T�%�4p�=�	��_
�B!�.�e:���rޗQ�ȏ/�/�h�U�����'�|�jG.���v,T����\����6o�m�	���G���i�D�2&���>�Q�f�7�O�λ��gU>�'��ȜF�b�KN+5�����Dy���e�_��W�j���C"��p�yt0 ��	��H��w�,��[]�@+G�N;V�a��Ew�#߷�|[�`]�;\����I�.p�,�x��T��z1&�� (�HGL"b�X�G��E
��+C������L�8x�qy
A��	^\��f~���}��Bb˽xA�������'p��d�/b������oL���mO+rIi���(2�Ko�ʍ;�@����N4�A�\��6����oeYO]�ų������R�FL���w#��Yrߵ8����H�p�k����(�W�