// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:16 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OG65RzBf9oby2SexpCy3N73bwQcE7lJkAsHcaXCvHusAwqrerB1TCtrqUsHTgK5O
zEqIr5zYdWCuB7Rd7Ol1Iv/ZI9WYttGYvNt9RRHLcD3knEwDIsK8iBlLL0aFsu3w
Jq6nQEzhYfu1e+QGZnR6y38tzfsbbf2ba8QFRa4aPqE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9088)
D6HAkaiQa5J2d9LPcQcvJMxEAgLMSnhqUUOCKWbU1CWaZQMtrtOPfxu513spJOxw
2KjCptV7CzXzGQkEVaMX+f5xHUM2QQdwwxe65Lxk6bJl1on1+dR6ncCiA3srrlOk
o3fn+QEpLqLwnrgtgAV3DJi8/PqlGs/gUZdz91qY+seI9vBjI+X7Q7uSniP4zA+N
skhah903vL5p2xS5+pYh+koWPJyUR52NsOUxbUEvz96qrYh6IOo5qFT/Yufc7nnu
zGUNtbhlQPBFx0Hi3RSE1xv5zbnWQLXmJyKdIx0HOzt+BLbMLxpXS46wLRwVFQo4
VEZ85iyc7mN4fBG32H3D7gHBuOJgU/XlaM0R7gY7ZG0c5Kpk04ScT6HtEO11A5Ef
oJ1luyl5PXe0ZJpsV4OITDcUGTeMe8lFeKx7j6K1otI+yBMf9CD9mu0Irrj3eeSs
WGweNhaP3ofnrAXPAydJhuO0DHrbBVzw3vm+T24EoqzH9waUTlRabPctXKacHRcQ
KKuBb2XBttA2JlgFtr2SD/NzMrT5PXmRSyhmPE2wg8W+9zjSg979pfv8PSiu60pU
g3EN1hg3/R1rdMOsAiqoWXVXyiIx4dVOihBq0in5x1KSKZiAWtsLUiQTPsMraoNZ
PxWo2ntc/KtepVKmgwYC89oIqLe7WQZ/RF33CAoadIe/CDmrI+AIryMBQ1hajM8b
sTtNCt+K0Smyt8ooCX0G15twj1U/+3ah91TTTJ5JC/1LH8gkOEU0ilizWuyp346Q
J8YHNXixP8pIPauJaQSBqOzg0R6NYJjVByD7c9CxOxhKe9FPIPMBm7O2heAbUWTN
DpgTdMMLFwCK34g3CagDBhv4uJcWwD+ULZgfbVem2TvjBC/qn49kiOzoE1V7rLIB
e/0IPBi8C8wOFGChauFHdk6Tb2q99++LAOMW8b+kLpk/a+Q6HHCzpG7plL3XH+KL
Xogz+cZuuZxgjPrEqtWd7t4ngSfGhpw1quft7DqPzpT4Y2FZ/T7vUG27P9fmq1Bo
OC1tdzGSH/4KN2VNd9cYXoe3W1aFZh6nex0loBulclIIx9gbHv/6N/ydXduoVN3O
QT21EAyeGmxOeijxxo6yoKfhn7PZTPWC+BBrp7/XPoCUR7v/rdR5P78qkrt8wyAy
VASxgkObgu/t/WuvIaTj7LZ8gq4IEw8lgpf+dMeCp2YyBGu8FA11TFWsXDTTv3FS
hGokz3Oa0LYRCM8hiFgmnq4yHibWCPHbaQB3pMpCsJuXwoCML/YwAL/XWTwjNyds
igcMlWe/gCozZSa2f/8pw0f7wiYhvyia9eITxYB+16DD96QxlW2itGP8YMaZZrFT
89szjDfDrYOl7ppmV9xSOK9fa1uedztYsueuDn4Ff78Nrmxj1B+de1aC1yvDYbCC
kgx6LHeC7yDHk2x72f3WTGeqnaHB4sGqXepcIZljmxVVs/HrzCLtBdidKDvsHjvV
UTtLtW4AF4OUL2XWBVVJGsRaSI+wWek3nI1WQchgiFYx1ANs8zT2rayiVsa7oiRO
6QWgZN0y27ywI0X/7EKfnIbTXVJHzm4bqfBdh6tRivkxa5vt9h0pcap0/z7LmNMg
stx3TecqAlfnS2Lid/yeqE/m2A1uKxTEw3EJuyjMCk0uhdlotPA5yU59rZbWdSa1
KFg17WO3Y0tut/z7Jxw25ksVz2a9Zy916hIWPV9KeAtRL97FsIQXtMGX4wgV7jh2
0mQhyADDqBiATmuu43EO9Ktw2EFdU4ZsV/ez7QXMji2xZcdXKZre7LB3fo5gmbOe
VgDDzzdS0lXH2jb7ELDnQfvlRISbcykx17dEbDlfgIFxIEHQcX6LiyJMpQYDq8xO
bYnDPNpdkgt2f+TdQAqlmur3jqLVWahFzY9Qv726gwV+ZgYzOkPnuCN0/ywA3/vi
uaTnTkcmOdX1R2fcRz6w3afy1zGQLSxdliLlmlRN762mKFNEwHeJ6mTJsXP8VomN
nlCCoSdVNd9ecN6ThML2+Q/dcZuxmsjizfCWVMmaCynkXwjpmuPZJztCsxivBN2a
5T4jCgW3WQrBFSB3Zl6THEqVlvdh1tSr2tFEdl6jPYLYiHw8RML/MVf/RaHwTrZZ
e9uO+CwOrPF/hYxQC8Rt7usyv7vrghS4O1a5fH4TFrIjDvy19baIQp/BuZkzRI3/
wkCoBqeqe0caPHu5yC7xvcecMzxfpDo2xC4pWA0r8h18vSaDiE8o4pRsGV9fZqTh
avgMEAwUaKZvvhJWuK3sYlYXQnGS0YO9RLKXSeati7+tnEQ5wWTKJlKeDZeJoQAX
cwTH2puJLQMnIpkbzjr6zCmDtMjLnZjSzzRMLaWGIuAKnk210wNpRiuIrTEKmucX
PX2g1rHqoW+zWyUMDlTmqdRNzPYzrVsRZsSwY2/tRPAwL9bDxM3occvgKOn07eWb
PEKcM1qOU3GjMoHz9S4bBtLuSOfe/2dAG6/dXhzWIxctAzFYBrZqM+KgCbsg1PoE
IjP7x+vpyYiZuTP3PjPKopnn+YTIi7Zk6LgawZ+uWWonj8TU3dxe1tFJGzX3jk7q
cOVSKOEnW9nwDlVz8+fH4G4D35Wix4TgQWX6Up8m559ShKto6FGX+cSF50OBSo8z
gZ8lnGsnBKrsBlYX+eL+cj6s19S9EMkTkE2IMCBsQLVY6V2eDGL6Fg6tF9BDr8gi
qhniWmh84WDqAHQUg94qaJPMeYZM1mH6jRCVhRRqJn0o5iSHxavbbCfOA20kgr33
roFD8xTFoXaYvzhMxFqdy++26kWVmEWTsUBgQ93AxnH959uJ6LIYvDA0MsE4EtJ3
KQvmJRermdCsnzd8kjV1Rbexy/c4amEs3lAnbqj7K8jxxb/fFD+9m16xDfzRGhO+
U5zbO/jOiMJyD558ieTxpmyRsoI7qyMne6VYDKKTaI8H3avwPHGE0KXY0axi/mX9
Q/H8F86vbi0/9xDgqYv47odxnL/OlX32r4+dcw+2gCGGW8Gs5zOgvzyTXyKDEzRJ
dGZGMDMrY9KeNJA1fJfkS/IFFSRqSBYJPuFoo4H9CbZZ/uNpYe6gcucV0fkT13EK
m507FwH9LzYkPzp2/cAeNh5KBJ9HR83wVt6eBPpMKBXRAKgDNyprGbOuWHqZHz8r
K63gb7kxMHDn7t94k+jX4tIzBbsq0y0+hUkUjA8xstVxw0heTKnjPa6Ntn41QgIa
pQgZTR/WVqH0Rw8T8Fy4gR83VqBW/qLJVgXv052+iIFIKdbORW8SwF3I+LzzQiJi
43OBsi9Jb4Df8RnnMdgAgU5PxNYJwvAN10ROHssSrwOjJgWlqXLqF878fAP3MbV+
29hzbTd6PdaVhXWd5wXXbyFHzO7h4DliyRK8bGH2V+V8dQHAaRrm/mB+PYMPtxCl
ILxdo2xXCqMIOKjXy/2KzA5+Vqx/Tba9t5VyiDZuqSoqYv0I57zhl6KAVToJHph9
/Ebff+RAQWyHQtgu2jFF/XLqQtiYJCtSxKpfuE1xsv5uXCS5EBHuU1Hp6PUHgxn5
4opkz3kzQP4A+ZQU8QJgllX/7IeEwKVpbWLHZLHPlzdgJS7E+m6TcHnHP9zCiBR+
sUv6m16ddNvfqixFR8klge9Uye02BmekkjPIHyfklQY3Guf1g69goZDQNQfCZhzM
9m6V9iE6IUay75Pf72JurOdDPtjtXXM3QpKV8ifxjDG6qziwcrujGY0hd2WCLn5j
mYqE6g9NF+Jh0Xdg4E52eLWi1zPpLscnDxjrxSm2oxBHXo1PHIBzPyCYHXY1ZM1P
QcKbKCpXWm0Mcd7chgCg6ju/cMFBIjdfYgyjbUHZGnW3v0Zm5+E8lzbqL5Jc736X
csYj6oZHV3X++TeLCh5D+RH9tCJ939WF+s2+gMJ+IT48ZCO/5NCvS1SJmB8QNrV6
mOFSPa444yCM78soa8jNTl5eegu072uI6gathqVPGMDjycKUhAqXb4niNysaWPKK
hyNgyfEtmS6WSFgBus0XfAoMzgnYtiQfwSp/vRJSff0xT4V7zYta2hJSTOo8+l0F
JZnfLasoYseclgUngbhW587NaQYh/gG4AQYTIeTOA2Xbqu9eOuYv9ONGB8RxN55n
YAqF37jgyPeEMav9GoBivBRNR7iikieqBdLC2GSk4FLw+5K3WO3IolGpkyxfSH61
DtHqeaMz5tN3pCPa9niapjbwwhjk7VaNbzLhB4EAlTLe2PDHCJPkC/85xvUcxfYC
U3IVN2hnJPnvfxSGKw+wpeV1YRcl8rG+bvtfKdedDaiQf2LI3DrbLMvUHb/QIGG/
KS3liSw92ZGhi4BsJKZaGYpJXRD/lCHnHKS6e+u98rZ1srYEo/EFS9BERjzi8YDT
FcxbSDqUFIt7tjVAaX+LETKEbKuavQ68g9gf0HbbFQLpXrLONFm3tzVQIfV4UAMW
sZibDqX9k1HmyWTP/ufOnSHWPwgjdUoJQVwiVKwcHRxsJltrxPJ4lugUHQvDUolU
BnIvBQTx6JbUDI/FFq7TdSY53V844UUmUOu9jUA2r9FExf3MGYlcYEsCzb1nMfbK
iEfWqbD4JeuIzaZltm7uZl9nyZtVTTziZIjVpVkAmeUmB6mMM3Y5r8vG0IkfcN/z
u41sKOka8UA27SphaxGhIRUeQ37C6p7EKEcm6jhQYDWdmb+4nwfa80SocgeuY8ho
BmQtcxmCuQVRhxo9lBf93wlYKrINDU3iIeV1p16ooEtfr/C57D4ovZKC66YeGC8x
9jagl6vm5n0f3s8CIoKwUK3G8A0IZfgW6CbIFY/ElPoB43+YC39uFWlYWlShucln
AfbfUQNkrbF1rwy+aeFAGbBhR7rb3EOPF1PV01I0OKH4CnvoyaxHKVfsJzpsA5c3
KpU6GKqralK/JKLFzZtedpjjQCm5zc1P7Ufcro8mzax3TXvai2UuMtj8cvuCOjNK
GTRkCooVik1oAIKwChhY7YZ90kJh0VPhR6fmf8/HrkQ8x1LUXAVDk4E/07FUfY4Y
jA9k5tWCoavqaMJ87aCc287CYPr9TQ90UcNPN37khhxgVSfT4UYqqodWgnUnHBtJ
6K/J6Ovxs8WnnKOI+SY2Xx6U9J3uBUFzCtDNdFzff+bHzAalWaCeoIORLy0yNWJn
RstLNFZJ1P/1QMe/nTOTRC2sXJuSBVjaE/BaTRynUmlCySIKCqimFPK92T7lbEN0
bVNWQ2RWEBoubA2e0Q48p/dbWeiR3rZrQmjXW1mnYG2YwZBR+05RO4vJGtRQDj8K
u+PNbLqZJn/8lxjxIenei1wW5jEAdkNIi4w2Mmt0+8WAUAu0VmsVerFTfTDFO4Ik
VlYxZSHbppgGlq+VlD+Qrd2DIrqZv9ezhE6Ru1ttxwuLR9+d4XLIXtvzD+vBGtp1
xdOEV3uj3QUvr3d1KnO1YfS53noGAw3vC3j91oyJLTHkWhDHU7UsdztCjyNjtC33
k6Qe4tcwGDfa+3VDAbMMuExqYTtu3xZU+B4ws7NpM8DwGJYzbELpF963pP8B9zaM
WWcYTKR+P1niTydyj8T53PYcHlPT8rWKtQo6u+bw6NxA2RJS9wYK3tCFuN+lI7jB
JMYb5UFnMw9wBEdr7pPZiZoxGyFQJ7BujBIjMjhh21SU8XDCMw70G1wDF2LTj8lt
Gsc1cxSU4d5VWRHA9lZ+SypZ6p9yRZ3zB9xQZAv+qTnFrb+inb3Gt2bCpZySQsj8
gJZdU35J6HKr/Psbev0V7KuVID95yReaBBDuqNhPPqbjE4Je8ER/ARn/gBLMmDBk
BLTrwHIXnwSofhT/xOS7+4b026cGa2ZfdR+wtoJEXYwbOv0dBoRp/4Opw7OtgsJ0
tEzVHhWurXf8FpaFf5gDZjhuj7OAd28towPvDhp7Wd3x3Ecd8T/yzAi2eXqVnZ1p
1SgiulmiqzIdNyO3xrcMKvUCRVy6GVngKXmxpZkoDY9CGP3ShBakkWaPbzokTW5/
+gPAry29Rb92ZToOAKg61pwrCu4w2+aYCbtxgOOuiJdLewvv4a2/S79BoyD/uItQ
2HfDEe808ElvhNGUDPMI4uBhBl2QDUukv5ssK+H1gZIgO0XDKIeYYufMO3cVvdeo
ncwo5UKyrJtg2WcWlBdxotQaMaTAECnCroUmGmcqc6BEEe86ORgBNLtHkwkEIpk1
8kDAaadz8Z7YKP3wkw/WB7m/qAXdf/wlJKlp7MLNMKxO0MkQ+yMMKIsFL7SLew8a
L5ShOnURk0/QB+pP37Z2AQLV39HuIkAFZrBtKFpm1seYWFBEYBgxjytD271duzwk
Wiu1aEkNq5s+e/hpAiySxFbM65OQ2zsvLxDtATBB/aYAYb+v9wSuG5cokEWRV50F
b6/oWuQHhXSb3dsNHAllhI61EKOXZOfdVrMnPgtVjNhFJKmOTJcwesQRH69GR5c3
TD9WftWZjSxt2sxA8gLY3UtT+M4gYfIdPFsghlyQIU0YApq7OxONk6YDSK1XY9Nf
b72k48IInIA9MxMHlENmP6H45WXc1sXW6K5L74ns3MccqDcWlmGH+GntRxmwsfvs
BgH4sl6PfV9hP3Tv+EAnJiXyFsoJ0tyA0R7AlNMuvj1RkYWkyniSIM1G6A+PXvaM
BwK1cK2hJLqOb9nl12Nkx8ZVmQ2TRw1X0+ld0fyC4HwCVdDJd5fgiLAF0ekLR3bw
Wmt9XRJSgKM/ee4MXBDXv7Fk4/CNAKMMSLV3opgk8PRJTrrzg8mk23BWbE824sf5
JeOSv7++FoyaY0qtBKDwiQfjvtoI0LFuLrhDfctue07ZDS+CczqtpOlO1bOsINxL
P1rf2Mk8xrpwpxpOrg+3wsAm4ytrLDt4oc+G6m3Aqs4WloBaQBoRu/TKD3IXBlAo
llxN6o5Ix4tcDoovXyWuAlaBamB3iEQfb3j0Nw0UHWdkcdTximQY+8FlvBgxMwGI
ShIf2loRw0dX4pnmySzTJUNXaBL7qbZadcvGGBaXnPxRfhNsCPLpYk97TrWY7rTj
V0S8u687smJsu1JSnMWJdD7kauT1s0w+0SKE9vNzxbSeDPQH2Dkfu4S9d0cZjLBx
E6s4q9DHEy1LifGrCgORMiFSsFVjS66b7khQ5UvZFR7LpOsVBtLufZD03gvoG16r
/qzuXV9HpJsr3dXhnP4tlAnj6RWHZbnviK8ybVmTwjP7RrU7A/8TDQ2+Mhc9htNz
YlAqrRaRgyT9IGWu8vpdxA2zAcvNOoDptYcXDAM5/oBDfH2TgZ6EW5elUrzd3Jqz
vDoujn9GDicIXkGOKGry54B9Y+D3uJww7e2DKUCk7p3EM0WU6u4PWBCaocNQ81Wq
Fc4XbGrdq1HtRc7JK6+GHfZoIOOxRVy0TbZ8NgRCFR2yr/AMEKBkqSoLRkrcukRa
ZHUUcOWSrNpwKq5K6hJVbacHqnU3FPkRLmDwNrAvYr6YWqkGqw7spEGqf1yNnQvU
X9Q9bxyvc0Ekgn7lukMWFa345lZTW716EmGaEfofqvMR9mkpB1wQIxGcgTy+1/oA
SjTyVmZiwv5zwv7rDiefZ7HJUivLKoRrCCtu5jvxsyXtTXN3pa85h+xA4L+27R1k
ovJnYe2kMyIfop5qgPsirj4jvcQxBzCb2mLzLL9DYJsrsCocbPpY3nSu1oWFfU8+
GoqPJ+h8NBUW/FjBg5ZOQEKHtOGD/Ug3I1XgoUTBrVVPcde6EHvBFkTPCE23mCIs
SqPOODk+hnnCj+ePrdSlZzCeLpB99AsLUppyBCENZPgVxVbjQnudJiRpu1yq1bP3
4Md493Xpx/snOyBa4JS07C4pmTc9qMb9jxsepeMPebmGCzu87EBklOG9WAomgcVd
QeNMQwE1s8bHTRevCeDO3iSj0wL/iSowg5O4CSoGkW3Q9niru6+3XVHIMVQxq04x
Ec2mKyyvGGjCLJ3fksgZJXYn2NJ+VZG3aGn6NOuj9pR+oDE19HdpVHHZZ44d8cIF
3MrIm3F05ZsOAC4HxHbk2gJ288f9RJLauO/KP8FdxFL7GO4/y2nU8zc+GaBmO/uL
lEaRIg6ups8eJwermR8fZoec0WXfT9Cn5YI003PGSTUCbv27lq45aCtg5hPDOhc2
8RJtXWfqSz580eVlSo1ulESiuVRcF+OZgTlHymDSuFwoCub1FekFHi9vdZIfSpVS
//YxsKSuuSH5+uJ3ZUX/MN4NDZV/OK6E2HG4ZoP1RoZO1VeaPlA5Fvk3fsOXEMEw
9MNiqN+Ltv58hj6levlES4LC3v44HwQSF1SKmah58Pz/4mU5KsGzfsawyhl5EExX
nJyvHekoWSiZXvjari7zix99u85R1ldWsIu5NknEMbf/RSn2aVXE+JbPxXfVNjgE
kLnBhFhbRbz9VrU9Xt4UJZU8r4CSLN6HDADhAYN1ypHWtZPhWYrqHxTvpXUySJLr
ak1YKrprCp8Jd5libBiYUP1brA9g06KhiPSn1RrcXWQB+n9qODY9WpSNBY+3hJau
IdD7B43BhuSgf9P0vuvmjkV2qgCC4ERhtKJUFOnoT/t9cghpqyaVEUPs7RTDg/sa
LvwJ3JV15+kdEDoaV5h7DVQmQYkDI3XiQCBzlFtqykBw55+knnfF23cjDCLgSJqr
RN5fUFN/QRUZlgwvA+48co+Ac0wVZ+jXQg0JtKRI/eX1NlH/m/2CIDgPMpP9+EQa
2emXkB6teIhd8duG+3FE1Glu6gihGyYArnMTovqisr+JElK/LPc+3kxRRWya+5F6
+rLNb95DbAVAZXaUXDrfHJJo+XzN6I/Yiig23a2KtcVqMWl4bZzbE14nj8tZmUYt
Kxf79Cka5gwsAD+FxIjrV7t+P1j2EgzYxPMd+Sj2wihGKlbmhbnjXWkUuvQUX7sx
4u+4MfGrLCEUW8+0r2jBzbIWFTKANh41WV+Kof9bRyQFirdvY7w1QyyXJnFTY4mU
SvgH9CA8LT7ZoCzfI+V5GQ0klJzSqG/5FDePigai1NPCRjEhMNz4yIYzFrC0HE9U
aUMHmVHsrkTz63a0QDqOwF+kmQEdmybVWTBx4HNv7Nr/HGWN0IingnqU13KysOgc
u7Fqg27mdoEnrA78utafDiu5rtnC71FZAOZtOfgZO5uPv9WkSuTG56aXhfZMt16G
BcWPaqgL9ISjra1vb6ptB8hMFVShBzlKc1qqDk8fxX6IlbYfcdqXgVR9b631H/Et
mYTC6cG39Z6J8eieXagsD7XW6Kt/g0xc8qrNCbOnbneSnSjydq7ufxyiN/xPwBBo
M8v5cB7xJK67PP+lyNYLrQROi/7PCCh0a1qLuxyhV2tn04YZvLD8WETCDvdCYqXc
n1iY20EeSwSAOMfA/z0P86jSQTMLHCHuHdGORHED9u/b26QMOC/wzI2HzXfRFwk9
8Z8RRtZwpjuQ59YUClqs5Hd3/HBp2C3tnnhZg5TkDMjb6LuxfO6KCDmIOhEjDFEK
OSHVlbCBocyrs1GvLKpa+AvUWAy9HJPH1p63wMHVw499+EyCeGtbvVc2pJEXLMw7
KlJ9qpg3Pf2WeCaOhWGUNFHgPahg3yogXAxusdUPD0y4kS7aiHGIXPlvnfCqCNAZ
Y6U2pJ52tpH3mpPsbVVq00MfrOhxu6oWDCnk5iAsDgbTxKft2xVOWF8CuNa/4QsA
edl/JCO4Ax0+HHLbTbzWhNbXUybhE94yAPZj0FIL2VQFQIJEaiRv1hnYvMJ7Dn1e
jWSR6CtV7B4IK6YjTQ+xDjgMJ18VJiRw/FQSaQ5KCmOc0dPdF9EVpGgQHO+eOOxP
E+pqsGfz6SOXxey894s/9KZHMv/797dkxRFobztpDMc3jeAlMJxzf+moZwWuO3w/
ZF0d97HNlsBOvZdYZozem9KYoyOSJU5z3hO9p30NBUjujqH8q+3c/eGo7x0mwdoD
yGkcCAlnKp1s4x3WmdquzbqBxcMcFVpBDXjsES/zjWWmF2mCEK+ONjRSqepRDJl6
h7aueM2Qz5/H1uwIPbrmOtv+rh95hXQ9zzFMKkHbILtx7u9CWaf0cbS9R/tGhoby
ihPDNhSY1+nFEvLxUb4W2OK4cHMQ8KhmWuKjhkU5yRxbbRBPgEu5P5tzWLWjapzR
RCvyBX0gFMD6n4/m9kjVmZP7pk8Gr9R9/MkmLpKqNcDb6wVy8D/szhTSyOuiJs2C
PDG6+seJ3mzGnq+Lsm73e3185C/Y7lGpeWWHvI7YOcTIUos49YpLG7fgYUGcnEbQ
L0sQusp6gm86BqMtE8OuWMDapSLfQos/goHJMmJrwegubdBxSHS9K6U+9X7dTxMl
0zDS7t/e4hp8/bIHz5OQzuXB1TPX4BBVT4q8QB64jqFbrwSxp4JZzoU7/vER5FE3
TgRvcwqEMKzT38dWtwQgM6VK80SO3EKYQMjFnYGkY/V0MA54bKwUurjtrwgV2KPt
bIqQGjItp6wRT3IawdjZEPu/6zDycZKOIu9/Np9MT3ARn40Zt+CMPd+szT9LDb/c
mMZGqqP2Sfdj1Ua5ELlhBwVDjwgvquUqhczgbcLS7WyBTieNCQo0rAJMK7+5LKpi
MCEahSYMx30a2pZLstU+TaDIz9GLXrNo0Qm1hcujHX4MfSXNMY0GZ5G4EINJyKeN
hUqo8tUfKEpqpS8RNgUhM767rv3Az+L4aHVkxiclfutkOvsBg13Ka0PXmZxciEO6
KNPcptroJQdwxkRcwn63agZqpW8vSbM/SrXzX8fVab5hMBpeVe77ivCVVwF63SEs
I+8T+1F0mFLcn3l0qahylLrIqhjn5UJLqZT/IGZu0G7u3/4SKbUWha+FY0uqg5NU
Ahb40PrzlHVZkn6w/Ne+heNTQwx9MctUT3+JKR61dV6OiN37vhwA/dPjK3K3I2Vs
7i3C6CZwqWGyW7FtuQugHgZRidDCcThbocr605+gV7xXWu0Z21wWi7T9MaBpL5Er
0IxjmIUegnD1RdqFcuLappq/3Bt1WgPYLcLHO04+zyNPtHAOQosbSKOmrLetP0xZ
A4gB1xouBOcUkWG4g/Tm3zsmZz6q7MceNc5PPSn5eMC3Dlr6qj222ymvwWyM7pMC
6pN/emGe+rLX6R8947ML4u3yNxojO+j7Z/1gHZeKBO42tn8RiT5xHm92fRjRPB9B
mCWZqglnhZRFaZuPamjzqhgJ8Cf7qyN30TK1AlX3AUTx1V2jj+aDHxueMpXYlSfX
Rp6VNVC2GNKjv/4BDj3mqbqwp0zETTFYSKBiSDwbr9QZWHxlYN7Ss8uwwRDQ7Tyz
3Ottr2+dQyNkBVBvC7QPE3EmSjSXAukUYAG9C3WzakxOU+Wr85yuENwlOVPSEFg1
4Rl/5WMu/4vD2F8DbGK9iojkAhUMBp4IyTh8xMT7rTOiTw8wR/KZZwTCNw6+FvNy
9iSCeEE6M8KNKI+glz+iuHez9goDzbsEOnDX3UGXaDprea7CAX+Dc9Jty6aR0+CY
RahZnHM6ETsUxzMjAJe7Xd3XLbDu1v46WJrQO2i2mFkRTYJS1S6cmTEW85sNqeEf
LoVPnWHp+BJ3tkVJMZU+Sa3dI0KylosdaPGmuRDatCY762lFe7TrtBYSLgJHtknK
96o/0P5kbusn4RWclP8nfPCtrfnv99ECYStjPsZE/oQkKTC2XwGApxVD+Svibko+
O0afausSQQZRnVG5x/6itdH5ICtvdbiPzAbpfofY2dCm95nvyCDXv/nCoXXm/Hbc
KBR/UGxwSO0kvei8XLndJX1GPTSbCcJJWGaEccp0yAKBtNGY6CIOS9DDuNZKa9MT
NEquph5TeTX+QE5znEnvhyrA3MizMEopksGCDl+D/OQDmHkN8AJZu5xGHMHlg+my
7pusB0+kZ2dTNmWxf5Jsc2pAO71woiIYpxhpOvPcMzCSXNGUOC1A3nhEyF96JxEb
8q3qjf6cjmCciXUlbc3f70zttuE+DcJLpdnXhGNqAH1MKn52mixh1QQxSNufpKoW
83jWlTnigvRLnfgeYv98USvqRSu2psYGvrfTEAbMcJrRm2dq9htCq0ZbB9ERR749
gRGqQVM/52V+zDR1Qvl16KATa4muIzmFSWS8kK66F3qCbkY70ECrY2rFBTeRSUQ6
Z84/y8VUNUVvcvSmj13XO+Qi/z4fNQqVCVfueAykGQ6Mv4tqyGfnWAySxHA7ftwc
bkctn5ilXJ/2qg+LqmHqkA==
`pragma protect end_protected
