-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
e5M/oW09Q1ivkwglST5Q6N/w765YUY4s2Y3uWEUzokJ8bwn4ic1ZVoUrPYskSitvuWrJAu4eK7jz
ID0eSUECLkgU0/xxCLHk87jhr+nw17Mn4r+q00KSvvP9QyWRYRtE0PWtEffm0sGIzlIqiFVoan0+
h2BLUD4Z4Yxfj8xnq91x2pnXFU95fNcpzKQLOoF2asfo5iIbnRc/yQcDt1Gt9ReH7v9rRSmctUrs
+cE1fSNmyElPmLviQ5AFSj8zHh74Dr4ZNoyNkJO+Rlezc+Wpdk68tX+NJDFyYZYIcEFFtQZCpIV+
pVmbn7YX+GYAxQkiyyi33fWLaUbkZlXnCOb/UA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8048)
`protect data_block
hGcxT7jvZ2vkAHzup+RlthykBg3tkVhyh5jOc2hlT/bHgeGQQ8eb1M3GriMMFfQGQhnuHO2AMFwD
iKhQ3ncme5YE46BvtRt6FCOguOA+FzyiQ28U5Qjjx+/FCKNmKKNlxWBVTfD10IXYI3AyrLWDAQ3n
2eBPaqHf0O9m/KRNGGkCJ+SiCIWPxEHUny4H31ssEWMw7zL5Js2zI4OCIC9D/jebydU34fgiiXbm
YjkGJTGReOgUGuOxn0KWRwxWbwR5OolOc2U5D63dlsKziOUDHJsPX8zitol6jo3qFAsghCWRS5bg
jvVQ4OCD3uu0jzl0an2q+UTW/KIdEjPipsjSJTeL5AdF+0yRBXSW2oncrnIkAc4+7KnQjzDvXaMl
Gab2tT8+ArDR9Vaaw8L+skr2PsI0sChCSScv21AfJVJ0seE0E8r4n23TUjeoMl09FeqkNqkCaNGD
a9SVS82+zFZfoMEeYcrVqOBq2SVdHcgXBuJ9Ia/XnzZ4POPfmqdBPxgRXyCkff46Z+LsnMhRTsBT
y7I+ebMF7Ib9w4AmRsyGdS9U3UCrj/wzYKNwwto4wv+PY6GCT5BOZ5UtyKIsnFSaMHrdwZTmgB00
ywHDldao+BtXxRDRHVU9XZcA/0Li5ipkcD/2E/mlwtfavvkUmZnm23yfdYykDUlfVTwnYEql8gcx
/bQFNkMfk3y1y0ousG6P91XEsSTsNL+HE8cKhrnhFN7pYxdzUmSqe1UQj1yUI/qwRi97z6t2mLi9
INisv1vMvEusiNwyyCHSf3WtTccHyP273sQwuwVztaWvMFR85DoYjdXUVhg//oCzSkY/c5q72Gve
KL9ZFFj0U2lQVxmsa03awN5k1/WI+thfnbCek1xVmPkIWjZ37aEgqyueIagiYQc6iNgvj2CNkELI
xSKWZYAmEZHlruu7msG83gzyqv08J1LTNSEJLnu15uLzENLE3S2pnWTlAd6B36Y+wmjHuoIk9MQh
dN3pptd+ZcbVTXdCoXdQre/FxbIS+qWW56tnC6JX9IMMV5MnKBE1Vh1cOAcAG5UojV99qwes0/lE
qcHAvVvvS0hwsGJWv+K4GYIyQUPfVWUFHfA0mxYi3FRKEc7y7M4eYHRq1bPFMY6sxofdYpw+4nV9
yZa2L/r2K6RLBKpci0DKTmwnHJBgclNHacC1+4mQliFaYiR16aYGceFlcp+EOBR6y87omURgY+AY
eYpxYqqfsXvPQy5D9oZ7GbfcrGYi5LNgs56lN59JpS0vbo08yi0+CJaTHk3mnj/KrIM9k8B+/7tv
dMA3sNUtT+2SDKL3SDHPTgqrIpN6dG6NzRA/MNyinlIgu3Y1Br3rxL8XLVR++e5zTHRfXMJREa9A
YfWdgr7jSWXwUWkihSOF3kxLIE5NOCTMtf7mp7e8PGKtgzPNkJtam99e/ASG0Fiht7iY08UFmEUc
lIEt0qTO9iJJFRBEySVlEjKgAtRaMzBsBBLNtSomheLvSIN5HOmokvOTsE8mnKefPzP6HhTJ8NdI
L1Z8gN9XChz2/uyp2vIOpKgaV6EqL3eW6FoOvqFs+g+DHje8Euh74WvS8HxqDRFC9cAU0KriQ4rH
TXxJFHW9wr3e31nx+b1A+rc20IrAkeb2RzoX6sMhm5ajZNiejYIXLAIrr8jP6sx5pyZjWqF8xq2W
vT/w6OQdRy1c6zKcidCd2Zcb39sLmoTLFd3QwCU94HCYdlv2K+aXltSY5CL8W2z1YwVEHuopKm0k
whSgLFeM1c9DNr6ujfctueztJzDwlq2mZUqhmCn/KQm2PrihzV5SFcNa4ejf/duGh+FS/8vyPl75
3cGkJKDyd7dTlrkq3jnvta49lO+Vc0282v1yu5zcIocqL5nDeLaSnsLfXcug+X9UCMXJlyLMPo8r
i6E20zIPzaRzVcjg6rqQ6Nln+is/km93I0mhH4VdkY85vUL+EL9NsU70Wl6nALruFN5ZrDqiXMOY
++HnbwV7DYtZ47H+nU2aAb3hOaDGCJ3wMB7ls8YAURRBQV6HoLOr7tLaekXGYh2JVV2LE0CF7cJY
Pj0eCpqess03IUJ1ZgL8T7CN6S5DgtQQb0IE+YMyHhmH62/eWaiMMCekXSfEcq4+UuOve2hkinJv
MjkJ72S2gFSNBS7d6edwMcxlj45mKNl6IbF2dYx3Yygia4kBOtUc4aejGy9OW5AvpG4FCkBsYI2w
mKWT9FcStlBVJqCA/M8lkVLnMRzkLy/ZRhuif1gQo0ED7s+0dk5hJ8SR1BvWk2K3p3Xkor94IgOp
qQdUdbj1PBl74+s3rbXlmD40B+pBDJo9albvh4C61qEX8PPKg/MzalelUOiO8xT1CFZOTyTtqi5O
sWWd+XVf/Rb1dTfjxg8i64FtTeeetpKaRtzkQMxjKOe8C9LFir/7yL/Slomk6tq64oViaIgRqepx
6CG/F3OAytsrvEB2EUmMV65+2avkoYL1lf2GgwV+TfsaKokFUOMo6rp7a+hAgx6QtX+lG2XUAiri
f/dJI69Hn+XpV35jWOzQpEp1Y/WlaYmec+zfoCWH1FfsBjNXjsd4W50cUmWTAwAbecCWXAknXvX9
81NbxgtmLWtCnTQKEE1GL59P7PPYJwsRHc4qfli6USs/iIxje95Q9oHKBPuNz2Jn9Qt+tN2awi3d
xyxs4kc9MyRqWbkSxFyTixuI30ok+euL/u5ec2pxBj8imobQ/s4qNsVoWg37SW+Xx2tVm6upr3zR
0LjgXbic2RWoSj6RNfSsyCMDKXqIhBc3LR0QykxroFehRn/AadpIYtkhx/Pb/R5qX6hu/6EVWtmB
8jRmPlOP/sCzA8MPhncNcD9ClAo7fBtuVt1SgJzAvIo1habrwmRQcFJVo2aBqioO4iEWSIgU1lP9
W2vS1341fqGTmvsUl4AqZWgfZRIt0Tx3EbopLn+JdArnnQk9fYgsne5aItaA+KqmYY7xBh3Fqa9Z
2WT+6QeFdWSHu/W6nRn1c3GI74yST8ZHhyHfzwZX5KJ1DviPgM+lVF5KMtUGI2iVbdk3WULxaBvA
kBXL9PPHL7Iqs7v/XqU722ydvKr6Y5TxCWVoGs5e7Y/R9KzrflibJlEJsUqXCg5JaVpViQMTjoiN
LyLOXH/e1s9GGWBFpA28YjMVZBYyvYb/j9lxWcAXNjWzSIhJ2IEWrC//JCiKnLpn2XToTw0cvmZ+
wAdVARK2zSvKsfyLIQ/Mp8a+yL1cAsLvjreeV3E8gHDawZGi/DLOTZAg7VlLW729yLJ75ahR7Ypt
5ZeaC/lMCr4S6WzYrSB2G4ySBD6RVYdCyEA89YvxSgqDnUUdIUia0PMozPa6YcIlyDPvKkLKI4Vb
ptQBWDyiPMT1C02Huznw9IBu61fH/ekVJUPqNAXaRedkVodlCKmpfsZBX0P2tS8a8MURZzpTphzH
rvjNVy9KNSpOkhY9RKPZQV9P9kqSZos55I2A2ELhG1F1SOmlKSyufN6bvxHCM68WaLVMBevyaHf8
YeENklXZ9UUliV33Xc8XaECXC4CbJ6Oz1Kr8Mohz8W3D+N3NGuOJHsO0E2JfuaYLddmyX0LValoO
ZkV2cgVSbD+0muRxeJ4iSAN5Yii/7ohv6yJBwMjdjQ1Yf42dKB8WryWcScgCS0GqyYYzxVjzlRZv
BUwWcWlGRoPW4U6fIi2m+/cActunlUJiSgfewfPmfzufOh6P+G75KF4NzPBi21M56ZRpjBPvq4A0
SZRniW+9leS5nvAVsiBJaoekN0jgbDROBxsI65IjEss9Sjj5CbVLjyxDDXitQEP7A8CgLRT+h5uH
bZcmTCSS8TrLHHZ6slS1Uogu0iMLz/84LYwQ/lV667IAZZhcSiabOyAK3Ljg4MqnabxjcOO6t4yx
h/9Vxn5vwEhZYLUs1IELrK+/ax9qD6MmJq+tHOjnkZSvVDwLU+Dz82Mq3PIoc019NgWLtWnfbPDb
8OWZQeoQi8iL+WFdCec7pnH8AIplcoDWoZYCrjoo1IjbWcX+90Ur7LqCrvWNZvWmGwz+U1pG4hPu
xSBR4zSmhISX+iwI8zYW6p9B1MwbHBOvBPjdw9/KdEfydi7mDXww7mWo/Zjh4FV/YlDZkcRttI6Z
vtig0n0/Arc8c4//fliffOMysBfzrSU/fkpctkC1ZDwYMJzT5Dxf/ojrSP5mdY+4jbPapGDvFVX0
O/I+k8CFNioN5XdiN0Hd8ciW1cAVxBpQ880HTX5IYYTbMR0h3y1YqhBSSl+1u5G1yFBOfLqhF4uz
558UTcj+mhUZu18F2sIDV/ggb9hcNZMZ+sM/n3BVHVv2ti+C/TJuVtwuAPWF6MSXjl9T/HnVUC3X
QBky81GFMDVL7btP48JHyrDFxZPm25H5h0cedNHiCKpFf3/R3VGvi2OqQvwl3izLXo5C3BbLhEzz
EYnyiyd/o1YBArM+xa8dejF+sm+Y3PnD0jBRWizn7CwUQLY8NKBlyQBTBe0C396I+tA9LUKfTcBU
rW0ymP7cmaV1rqOsZKIemTomgw57Bj/G1nZlspyIcODDNTVCoBf2j6Bgw7hqzexYyN/XMEzhI0E7
8keXExFyQD68Nt21/6Efxl0JcjlfPA5LOKfX3uA2xNHaejLQyPyacOAtzowyHAKAfPtlGNquDqbA
SA/S53gZgykcRsIU7VoNAepm9GJLb4dCCFEXF42VlkLK4M5eNopak9p5fw//Q03UPPzH+sWLgWCr
9HZcD4VUlVOH+CxZEIOzu6o95+HpUkhLZsPsBakPPiYF6s3EgMjBenGL2g2Y8vG00M7g74s2tl8E
YChcFAYwSE7PQXEt4Yy28NR4VQ2eGvb/wtkL5x9abPpsBBN8/v9KTLwqyYCiAle2zbz+U4a/xjwk
BdhgWfH/QHiaYniyisMhWpSMUk4OnAHufmjhkF3MeAe85056TKuhJl9FGu69dFqU3+PbkFg+7BDv
I5QygDYQ1/ssav4zv6i/k0xxjpFcPkbKhUDhcHCXCGbVnisqD1hMMPEyHoAOQAW0AtesaE/66mUP
jnhfTRBig9U3jMeXsKAODj1Lwsli2BKxTe+5nIzis6tUONU/40xD67+LfFsU2Glw++b7tQ0274h4
FVqYgp6SFdhwrVWA21ZhIw7Dz8FhxmBAdnZC0yhYNZHVXOTHwhUPkRHG/6KhlxGGpAJ6Qh383lAf
Ajp1cnMKz6zdmMbWz0Cl1fqNK2TydUAU6/5Rt0NJrjWegIUX72nQaJkfAe8EOYkPMNdSFdbxggLd
ZmysUZ1FZeGKx2cr6gVVpigTGDPBU+ZQ2jqtObAbk8CpbX0+utffaqUt0/i0xInxLayBT6RRpqRc
q7jEPG5zGEXztmchvDOQu+PyPpxWDXJiYBgORYL4n+g4d3Uo0A8gfzwBZv25s06BOUS5xq+vjr8n
u8KC0nYeqlK3VAZeMxwlzKN7G7n+0nhxJZPllo3Zp2YeopQJ4+UY86XXrSNa350JLjIo+7P3FmfY
LBQ81RFhrz2fMPFFfZefd6BkJMM4vy1Z3c3Y2ADii1UWDNxOn31I0vqKRaZ6ryS4HT9wZIBUJ8nl
kQQbc54Roj5wteLdGDOP82YEcjUlepK1rzCPxPgnkGZBA48cjz2dB+KGS+V+9rNFQ9T1FSq49nJ9
lHZ9JRMwNKoOMCC1NIfiZYEImPjyR849PeAzNXiy/jyQVoLvPDE0WJ30qpGXweNoByWRph0xDTqO
IaRqbexjzjuutJmZii2ZwNLHjOPkKumJ/f6L4G9tWTZH9xXCaoQhjHVvIofjyc0G6EiKaC2DTaLF
5iDXJEksnhnGS17VAYoOyNBo33VqgyYb0rpzQyhEv+FZtDfFYZjbunKv7rXT3C3H6PKDDq2S93kF
Yzvg3tjaZaEv6lWhuBUZxSdeJGsuYSvj3iwb6E1pluEp1oogDTNIdjTjGv1cv+HHV0ZUVzSdujIV
mEEs4qYU0E92glRMgH3vBtJpB7K7nabIMZrRxhbp6Icy4BlybTOo+gM5vPdwGXS3Bwy7/elNINme
SbHNzH0F17pMkAhtoXkp+Vgp5pTYZI2EVeC+Gx2uWAG1QLIP98nXxrYJQLpRB7ejJN8wFtbhnwTi
Jw8XBybIUwpS+SqIPcf/SjoGm7LMEVWqCJd7nh7QE4/xOZGaDSNpjSg7rRdGYCkUD03sTJjHfZGQ
BwNMHXmw8O5TdUaHbRY8AVr8M5bw9iJZcePcIEjYf4NJRFMML3Ma6qU2pmF0fJIPYxxCuFQN+4mM
43EKgFzKGJ2U4q1jpIgJriIlSSjkKmNTGUJyYwPD2UG7kqPhZdaHdx7yAoT5DzM1iRp9cep0tbC4
wwI8G0NszfDvN3ayQIYfuwtWLirsJu8zUVc/8y/A0rfY54Mt69pJUQZlzTpEtpvza3LA6LkmZv/S
SuSUdXWpxOf61k8vdrKL0Yrodt0uzHtfcKNvgL0rXZ6cnCja98XjWpqGTaeIKrRsfkioGe4zDsaI
Z6FZ44fkwXqk4+PaYE0gfdTAZaX9Bc2qpPs0J6U1MSlTCqhet2Ol3t5B/gOhIw31oz8vmo/8rGhb
uwaMrBnz33s0zot0dkk0BP8D73y8MxvooQ4Od8whh6dvIK+v8L2wxuVCL10QWbl78zLw6rnESXMZ
6IbIlcV5UwA+6rZXKUdTzpru0m7YuK4VWWu7nsClbtOLOkmeNZF0m/K3Rq3oS6bTlzFvU+nlHzVR
amO97pc7OphJGk+/J6kE2tA/gqCqzEUTzi2al14lFCCiTVIv5CoHVv7LxeLgDl5sRNeUpvddVmPX
oVTzT+14UB9CdpqXbfVrmC2p0/IMUiPZ333uNAVYdbG8N6MCXR+7qO7uOLbhAeJOk7iyjWVmCOFV
iIQ5j5y1nhkGxdh/nE9bjlHBz+aA+ShseAQ3lZwPlNrwVqsI1Bl0PKw8o/OdBPjTLWCyLobHtBnl
0GijLVMAhTBNU7IkrFvQRWQT3lqkfUooljFij6NGsPVjB1bLKcJU9aY822reUivgNDzFCor8tP2i
2uzqPwsj/uxVl0odfapKJCrtkqwWTPqwt7uCaeyUYeeAO13mDHA4lgvvh2s1YqCA14mS0g0IBgSW
i7viy4jzNeoqODYS3k0CX5NluO3LUXigutiW6v4dcdboHrRD2Awt9/p2YzRoFglw7DgLuaxLk/Pa
Bxh1ZVT+mr0zG07CQQIpydq+9yiapUe5aOAUY6+5v3CzHrvEYNpOhloRg9vu4nerINofAG2s+zB4
+Eg3SAnV45WYphFDsldYx1j8SliStUsvoWoQ0F9vgjaB+phdHY2W4UwB8WoPEWJK/gBnQa/Eywi8
CQNx2pyhYHzXxdb9LaKHowQcik0NW+JMwWz37aGoLd7ALeCIRwl7KT/HWmj9mI95cfenfPpz8rqp
V70yDDPQUklmm3am3iAy2ISpLZNS3Jnz//TefSAZcCrPHVD6N1M1zMPsCX1UqNNWbWE+p2aXQeo5
kB+fywspZNI6FxFanlMPlKTJTbMZepd4vpuUJQVE1U1V3JCp/ibUc4J10eBY/UkQsGWFvyGXa40S
Qh9rvRaiHYs2tmxY9xHQY1GV5Pho94Y+XPu6Q0QfIjzs9IVHk6s75hDpXdQxLDw9bYmom9uQF84s
2k5OpUgrEIrYJ5nfdbcKmimT4qXecQu1NK1eRyE4WtJmNV3lNQZP2ppF8IPQZOeo3ddaqq29ERsO
WFh79zQZ911nfCGqG+nLYeXpYsG2Pkhog/DdRNVZnYeYFUH7a51gUNYkfFOACtu9uAMkuXjiz53U
Ql80xoSz+LvvibKX6bQds7PohTlVV4SPrDJbCw+kg0f37Z3OHIEvK61wAE6yeJupGqtlgSSByD7G
n1O3Gu78001kE2SWerrFWUGWX1PhVvjm94vzq2QXPayrPP/mhO+K6fQ3vTvN4JuyelP9AT9B04YS
j8NDjQVPLfoXU6/C6Tt0Pq3TV71Eq3yPR2jP68FMPfRvTnRnzNeIxGJtg5xEl1DJK1KvQXwv7ykX
boTb4oLDOXXzqq9kqkYK9zTuS8YeDBKmJweQ1gNNQlJCSsApCl5miIrseunr5UQJrEjug4+jc9Nr
RTphxTDRy6284Mqrs2UEwXJeKSl/yzJiCYyy3cFeiORogfuyUT0qX3dNr/J7X2zpRpVDvDDIWfea
6wVlvK8/fAXx9TZykUruoMtcCMUDelrHKWaTp0lJboVv3sqT5vL7qZzLaMQYdYmEJFeVp9Pxd/po
RmcaMJ9CPpdalK2qQU9mLs8Q+Ot7rTz/AnCFzBNV6bKriqXPUD0fUSLboxDFvtuQjJpcIQxvnpSV
tJwd2QrL3apfvcmKykjV71RVqgL6O6Yh/Gvzip1bXv8hz98yC7DmViB5s/EGjwBkw7iHv3H3Zubk
Wz2pORDuH43IwLf02yUgKC5HCGOfr5g6jGGHhImHQWkiNgYnOo4r29+KkhVx6kduDLXkLj1oe4wn
8eKl7KBweATv+/UXzMbKt5ycgTs23Lk2+7oawQf99kZJ+PsUlA6oWxMDecIvqQuMQwPlB3wrQk7n
Al/R4zR5hAVI3oXJIsX/fyda3xDKyHR+s4SWpKVI1yLb1QYFtbIgLZazQ1GUOjT7iMfnXoyooU1e
xzW4hAUJEMosk8xY3daZkAucsG51yRmdZGjRJzkxh8TSkCKwCcteJmQIBIozWr0I8OE5rGXJcee+
BOg16zhzTmlx9sK22EwQQ0zrQvkki8ZGcLXnsPajRVDzcmHaT2g3ET1UzpovmBQlm7pB3ejRm2Ud
7iD7UHBaD3RwQWhGG7BCJanNMDRCvN5O0+SGpkJLcupUG7B+VKhinRTDmJk/P74Y6FdMuU8c62xx
lGF/0kEXRo5UNsAswhYThtwAUHPhfertKu2JVDPCAm7JixgksG2DI74FSDZeu9Y7wAfZcaKKI0f9
X1dImXZvbKxP3Tqav1lKKIIVj6rdz1ecOFamkWz44FPEZkIxKahSk0HEWkfRbJBE/WFK+EJL0luh
fopIS/1wsVSG2ON5hBNBPF6QgTP1O4ngbpfYVF0CZHDioNBx+27LsBEeyNZykIovCsKScW/q2Cqg
jA9h1Gm1VtFu4/SzjQfgvmMUZrdabRZxw8xzD0R+OKyeONGnRA0zuBwJOb0MzxQSAxdjPCc5U7mO
lgC+HCw3pvDRWxy7wZPbvr9RA4kHKtpx02psyMxND4pIFEPOEt1GY5gkpb4T9oMLOSaMzBJhcSs5
/VTlKDEMPy4QTr7CKglBeMdTO6Muh7FfFL2xRyNafGiQuR8YODEFELXgZp+GK+p3IICKcIpkTXpj
0d5xCb78cvgsd2yjliLJOcWOmx/VRDa5B/hUt+D//opmQhx2sbJ59HUWoAXha4xr0AtKqDTiTFmY
h1YQ420ugKOOlLb4IGk1Jex9aLJID9L/Q39RS5OnvT/B4fQsVdDdqkKi5fMljZcJJO5UP4hnf0cb
nVQ6B8w/41qh2MKV/a1mwi/Bw4pN+6R8DYU4T4n+ZihI0i03/7CvK6skZYWkHH2BNoUKxAHA29VQ
DT018Do9jr2qLDfw8EeuV7OOr8yGbi5Cp3lWIHpKZ9jRyHxQakTS+slyGGmdgPtO7BaiNSdD+1Kc
w/CU1GXUpupvq0tqe6DjSryPACAeAxxR5keRVE1lBefaGSYav5ZBzLpBcQiQ6/wna1mCcChtlXE3
l7y0J3fotRSQEfZSIgT8BAGx7RevQO3wSuUH12FGTirscP8BPD4uk7d/XQjZpGNfVK7IzZ6YtOwm
fksciqkSgcVBDljUA6n49BHzx5KvA42uop7d0NLW/SU+p8H0XjLCO7S78hlcpaivEaT2yC5mtZK9
MIuNlbx0gPFT/VdXLghyPaR0hq1s+Dz0HPZQIyuJfH9bpVpzWvBS0M3vXpZnfM9yetGGuU1jcNW5
HTAUAsqi2g7mjmwqNskxHh0jTl8dYAVOXeaul7K7YWyujv843cEqDuCZQXiBYbi6rdSqWIplpcr4
+Pe8KFfsQetPRBx52F/JATwQG+1UN8OohAxF361Wkt6BRSNjUkk+FVpcF9ZAZpdSay7fJyfEMTvq
B3o2dOjBq4g3wgYxHz89Cw2BEIPyI9NpX5omCX0qUjxNLyJQOqMFVxG8rkhQUc8W26GoX+497i+W
yqSUR7uYDk/i2PukZ50r076kabBgnLDND+WePeiJ9JEfCCw8evBxgzsSxATBi72lZT8yvf5I9jry
ugYlKF2RDweDZpUv4L2Av9qkMzXP5cp7CqB9oGPaauqei6CnPzDpYpyzh4ELnNkB0AyLxSyOvVFY
amaIGEsJjUwfORojhYNr9tublAiAeGs9RAkNIkrFAwAbA2sNDlwAqX5EiEIWSPOI81oLJo4w7mos
4SYwpj4GEyK175a0ReRq4KLEoyRxpk3BLGsOl0qQ7+3MC0k78Rz1nxhUhaZsadSOfT6mDN/Eeer6
RU28Ucbz4FwcQfdWkbF7b9AYoWFPNR56O4QT+4TM6yGaPKVxF/U10Y3iRPU4iL6d4adAeVh3jJay
E7KlhA1cwLHSpdUPp5QbWQ/DBJDa7wzFa+TkSypNeID4wtUniwxBqfMEx1Dn8LFp+vF2SXNWMJM7
S+GwVH1tpe+2D7jK02AuuTJVvYl9jlAreiLJ3nCE6VQ08PgENeGkLTqnvzQIin+mn1s3cilioojv
SQ0WhivlI5cqQdWeg2JJXeog8/r3b6X3/qLzGwRHKUE3m6SI4MOWwAhP2+tzOTsD6TrvrFxPf1PO
koxVhJjCGsjTriM=
`protect end_protected
