// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:15 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
on9DqLgc3uwDqVBmX+armp0BYoctLtucv11IfXWUuTMzq1J9XrXGtxytv5K6kFKo
t50aimxgL1CTidRbVp8qh8mLjoLj2tRR22sEzxXTlSk0Gj+GG+Rkl3+YmM3BUGRl
I/HKIvVDQ3unqEjpUb5NKwerqM3j42cHvfmkMGfNBb0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24512)
mztKz7QfzFODjhnTizvQwtOO63fCIMYZDPus+uFn3ufXmf3vzKcqM69n9nV/xQWC
t/dKHTTRft7hsaU9Gtpsajk6NEFjgWlaExDg5Wx6wVEmyPcmF5Dz/EqxiReHc08h
I1xfs5Tlcnk480XquEoRch0DWXLAWN4WT0GPNcgIzLKLy2Np7xczK2foBouniG/O
0QYN5itODSLWHSXHENhSUn84CMctxRENWOxDDh4qiVCMME6D5Ep/XzKlr6OkWRtk
hN4C7NXxS/FU+iNmh3zDelGHFK0r+iSWPK8NpwMT1zWXuoLVii4fNRfkjX2kk7Nm
N9mGmB9kstjFYeljmvTSDUCNjj1SI1UutIq2z/8jvW6PQQbyJMZ4l7NMVqDAv66+
YUwJrJT8LFfOLIQiSV8z8TG+WMCHYKg0CKb14r2VdkvvlytNlzvPL4j17PeMag74
k035pGWc/CGgJZgvSeWVGFtcwY99ZQXZwBAaybwcNIFhFiNZ7T3qR2SWK8VJ4mPm
HtOInycVMkb8ABeGG0NyTBb6e4FiD8V5xDmRA53Yo//cTT83kfJpkbxNpwXr0EKT
meMNLDY8meNx82bvCOYG4tH6G+Tc7V3drwXDomXZ1jw1R9+VUvCCjMm+r1UeaNy5
X6K3LNX1Ho9ZGUz3Azj7HRdmFhjNrDfCx5Plej5Xr4MwmTi7vgxCxMOC/h2glXrJ
IzuVU8RKjp2RtcHBH9X+2eTQaJECNmsi1s4HeoEOu764+XxZEzlXxo2TFMvItqIN
pJl622kVhMzSe26q3aFDnpwjQNZIVDDt/lALEF/GFutpMaIWO6APfh9OleC+m6x8
SY6ABU9JH1OSlCYnxUvl1M3H1OJekKAESyE8RLvj/bezVKmPOjpPAXLGLeqaj/xg
hBsXLwZwDFOh+YUokNyO91z6Z8ygYefW0OlWGqqvYk0xVlqKOVLGbYkCYGIe+6iK
ClHvTnxrePkgiZgwE6aLtqE3cmqzMZ3DN5bpofS55LD1+9qeolrlQWtWrCgFDN37
a5HC2Mo+rZDG5l6RaG9gPZXScERn3lVbzfMQCpTNexvcv2G/PGrlosFrQUUv471M
iIJxfQvpDc6UYJOull4yGQdklgYF6yNh3EP+/1WolfFUv7Dr0vT4nPsd9gr+fLvH
3wcF92jSI4ghaW4ZmftEVQhXt5JGD8cFklxyHnuemyoq80NJwfk/87zb8JkIcKnS
lk1hdRndaNbh3/U513Emykf8hsNZuvRMiXQWqrQU8BOXC7u2mtNM1YlWteSd/v8H
qSKGEAFitWPbtdS8oyaKC4Bzf2Vjx10KF/5jWEudMnzedbnZMfzk0KMegk6ss7F8
25whn402Z6LK3fDp9MxaAqWweEmBd9KHBd1atMAjm/nHpPbPlTCA0Ll4izueQNcW
PEGLqq1w1Y4UGwystC67HznXDRtWh/ZBPL+KmifcaUetZ79v4lbWnGsy8ej/lbQI
ZSQZL43U61uCK/KdECiLzcabFsAOliPE9yg/dnbpGRIeb2VJ/1SicYIuAiFJ0nAY
SATuaMNYGuuKfRD0DaGlfekN+YLg060gcUm6COk+wcHxE/kFP/9f/LIUP1ZCRb5M
QP2poDUZLJv3K57rqxvJgPWazab2YdwDf2wyMvAFSCglXWzQzhfWvtz4bNYWkXw2
q4pigGLTUL7qPhYtgyZgF/jeAmfx9GmDVx1ubeDwDReP15qLNOtMzS2qShoMr6HM
qkySmbm3aXrm38kClVoE4HP3LagSsvipPQpy1EcTyrpqte454qVRFFonFWJSioDy
MFcIZZx78uLlWlXfjgnv1NzKNWUpUHxEj4csfMgS5qtrkFRaXy79cHDK1Xb7CW9X
uLu8Q16oO7oC9JPqJN4WZsU3NslkmK9RaIkZ6VHcA5mAeeYX6PhnPNeG46FEedvu
bcYP2RLOPeZh8clw3A1adVx6lQwpsxC23O+bN6SE1a157rBzKmHf4tPF6LHryegI
IHMB3Rlyqb79MTbiD5QBGq0Z27tRIM9//sxa5rF8Ls0ODD/0HwmL8f/lcpF4guz3
U+GTojoZvnq3SpSk7V9Rp5XCpZRfFJaYgFsEfEBFHYMX7m/cBGYkKNgUErnM2jCM
9DRmrT1pXjX9drhODgkvqoZhwMsf4QSp2MTufiVNRvVqM8pm+yFIyEyf59b3e69e
XxEVYziP/+iz20JwoxRGvMF4KjpICGjEKijJqiEIrCgl8mqwVXDCXY9EIUyfNjR9
+LIPtDNU9NDChRUyDGYE+oKpGm4td3+0pGAWoNwF8vTGlBJZoNAaIxq0oWSPOiJg
0UvX+POfaW9qn+UYSxJDQy19ZNC1HSGmcVMFRszS9SOlgUlX4OHPoofKGWWxvytY
fTpumGuF9vWtnlX5FZhWb0lRQzFWB6loX/XSyqd8/gjVELI/P74rf4KAgv59GLbm
fahlLN48EvZt6sU6bFEVQUL/bBRJLW6RyG//t2i4UJzL/sc96GRCNlySs87YjwL2
BekdMl5ll4XOjuwvRkGg+WNSnzz/VpDqavzbUHuJlXZnvZOGDegK2Wm5B08/1xdG
IgQcQ7amtCml5laa7l8JPElgrqd/5quwPoscQpLoUR8n3Zxqg9fqkgmEbGVNTcsf
7T2n9hEqG+LRF0IvXBmnLUxoCurR9woyiUWqpSN6UMfd08KUSdxXfejSc9Asg+RO
Vg8+WYuX95NEKrdcCAu+aYKk4xPcuoHaMU/lbTBmIRUUQIrQ3Izac+F6ZG2pA1d3
nIhwY0067LfSpC95EnU62uX5ArpQTFqL5C42f0S05fGsKhl0RsM+GhVLit2EyQmA
IEUBTzg+UdbgeZvgYP6VnudSo8PTXUBNPV54b5sIjzVwRQhUfzOZ8HiTYgK3PEHF
+G2kt5OCxhqMb6ZEUwvg4wE8fO6j/XrRxQXX17ETucya5yPD+jRGchQMQEJE++IO
V8tHJtvNa/RQQ4u/mKtd0BTQbZKZQFpzfKARfsKerU6jgB/1iFmBPN/rFortyJVA
09+uWS171vk5QlGln9TKQvCclGgRyH7KdA2GueqOJMukEcnzpbiO62xYvnhhFcA5
j2Jv5SU6w29AZ2v3/RAVbgBkoOV7TUH0sYN86e5U+jjK9GOjv1xBF6dTDZuM+/ng
BRNUKYryraVupWHJeM+0fceyuuZRsdhdr2Wij9njWttepeOgcurATNpdKEYPSDum
zAs+gDbqBseu6kpkeDrIkK+FYF3bmb6/S+A2Y8AocfxfQqwLm33wotZLBBlVKRsC
WP5mJAQYmSJsRrDYyh1Az9smHweKgqpaK78u9j/0DaSKrn4HJGF2FU2s4D6TsFwd
lJq+41zKENqdAHyWkhfS32HbeSh6vQj5MecxXKB8VTQjJGtfo+ZKpbVtMndNsQ/p
Q8GXgsAtrjEWYqswnE2M6AZUQhUahe+1QUO2LeKEjfESvFCDycTH0UIagrFW8dSA
WkGMOUvHG5inQ74F3BXObHhwsXccjERa+VCp/G5DzSmYS7l90/0Uwh9OYT1xy18r
6SGxC29fNeCU+rEnCKhS93cN/zXrnP8vNGafc7IWwXu1Zqe1cpYUrbKJa4IwLcA5
6xSvMkMYGL8rZkQaiaEiqF3x0aKFv9XOEWShXt6/heiAC4WDbzUD4LZ2b+ysr7d7
GDrrWfSfcO9X+/WQmkKf5zmfFUvc3tA3mgMCps2LRlzLBS3gRVFQK37gMQJ5p74i
RDxndlMzMt9KphSIh5fuH03R5BMpUabWt0Pwu3gMv68kNctdwnOHhLvab1cjmGpq
VjGyFp5ATtknT/o/Y/VAfOqatFxTcul7yp6o25ZvFlNXQDn2ooFv4nAyN7RyiZPa
R4DKPORvVDZhSFMl7bZIcPaelgzo4ywDEEm5iqSYSTVatdUhdTg9fH7M3XEJuJws
B7qr/s7JlfriXduUBy4mdrQtNMdgBP5todkaklk4WD+LTGR6309As4W1h+YnmHUQ
UO3Q7RxOqizWOo2PTF7R9jNJ5Qa3OZKAKUeFWzfLbU/s/S1tTAvDurxPXg6rm9/j
W1CmMpMzqX7hXJcBYvbIa+dVbJnfn2hY2NQL8s+i4/w6ikiA0zI8P8S2m2N7gRt5
AnOdW8x+FKGPm/CCY86GM+LybcUr/29MQthFz38pqfK/Jqiimm8AtnsWiZ2MLJ6D
VLdGr5T/wOeZ84naSDSUik1huo4CfMMU9y5IkUuh8hOst7Fry9Ed+VnZQqLktSHJ
S2vzguDqyt49MemToy1qdCiCOK6Y9lvDyWMIL2yaVYCOoCRo/U+OH/DNxYM9TuQd
nSnRV9p36h3jHN4CKOtfLX1Kgpz7w8S24ngAcVVTDfNl9AWQPbzC5VNYuoqcmihT
3YlQAwYln/sUFF4lFYJpAM2Q+4jPBKfzTaARxjZTbBY4ypxIADSV+WK83wd738rn
EU0xo25iq3wd0BUoTXmfQJWna2PSVF8HmM1M2Yz/sivptZmwlpTbEtKfi+lKYJji
nUZ73FIXjA6eWRL2gof3YgWyHK9Sr8A2QqjXBIyhQyaO62wZ2nc4tP52sQdWA0Hj
+ZFiMGa+ewcYvseGTxhAq3Rd+io8KYrA0+BqitN7Um9UG17KPLWidWwTjF9Un11g
Yz0cl+PsysbegIkHp2m5qgnFy2LUtgSF3+lC8f6KskUyRpwOabqsWQo5bF0j7EwV
zBBGQGBmDaSibPG66vxzt2JlAErBwtao0Mr/5EhzUH/1Kq/gu8gdYpFSKR0ESa7b
mHf21YZ5LAUOmxH1cAuh2q3p6lijuzPvloNmy9cgOWQgujtzhpKMCTLemwBMr/NK
tRT+HtFrIjqFa/oxnOr3o4wImMGxoGyW0lGPhdAwRd4p9QjCvutje56WFMSzVBtU
+fbTwM/VOxI468tZNHPANgPWjwbSQ6W7BkKmwzQS24Sp4qhh6hOue9wItwRVggI6
cX+Z+zjxs/LRNdxiTkjKCK8Nr/BLPEQtA5fR3C7X3y6S2HsPp5xWkSUD/OMba+ae
6AiKEPv1R0MvxcqT/7PvBfiCZgzdNLSF4hVvehqyhbWuXyzt6kAAbMIKNmIwhh77
Z8mM+NhW51ZG6WiMS/0UCJNaPzASqEJtgoZWVW831ZQAzttT0Ye0vvnE/NQ8vmr3
hJQzRALLJ9sbdGQQvkOkNCHs+qga6JW/dywmVO2lUtAxXAAmHzQBjdArt6RhwHus
WOwYKtjXRM7Zuke+wjYbpbzGBQDA7ZIewD4IMdKWdyI4HuOt1OcwZXkPaXYZJir6
uReaKndFPMnLAq1O0mQmysUO4sxuYXOwP20VJjB1T51J0MsnBt52j9ThE2VTdCGU
dMu+BHq6ay2QRZpxFGShrg1x0Jl61XIT0wupYfwoCPZtF8Ds4tUH4B13gKbRMoP3
CNT/Cxir39TeQbSsiYaUODC8h5QstgWwU26wYzJGXtuVfYMDGC5EVkpF4m5HWncB
Cq3Lo3RfvUT4u3oRbKM916RZlcH7Ka8u+I7IYF355Qg8fd7Vmy8AlG9ZcAKD4Amj
spWBdy7vJLU5JFzw27g2ssndwJW3wuFmGrgE6qCB8FmECBV0ztMqVARrCUC34Afo
kxdNckK6cm+mPBZ1qwHTJL83dBeaF/gtlbPUHHe5nt73TWYAxIFQvEWU6vqRnuui
oYMi/YuGYPNd9QI+FXwMulxBuHGUC6raOMXs0vloIBgMAgKBmt/q3KLOpkETyXSI
NnZpiRGSSy4MgTjHEt+3TffF0RXowkF5ADgPjNxUsGrSpgBQOLq8GMN/IO8YfBrR
+Wuv9t/xxsCd68yp49PY+ek995Xq0nNUGznA2ClUf6BCoLhQGlKA/ZOAcCEfNaK1
qKu/fVGx2mI/Rqj7+HK4bkgNcQ/W0/W/d1jV5gO5uzvmIE/D2H964jGk+jIIJJrF
Hz7Cmy3OVEU0zzLTZEZByG9ZEF17dCR+5L9lLDGo6+3B3jLw3o5/0X7W6UNwERQg
shrF1ceTCmG7c8nAHMI0aAGDw3MPrhw0HFY0POwcaqc8iMLfA+trrGk590MHBCfP
/Vw54As1U90i7BTM9fYKd2CMnbmNv4SNYrweHz1aCMNUF0lglgt+aA6Xc33tLLni
87A4eCqxiFEHatVnG2Wwpf+NqlngkPIrl7FBZy4N1LB2X5QmQ5nyihtEd8H62qjb
XlUDrrZfG5TuvKhyI+MuYDllsEh3tdMTr2uN5BQoGqJ0+vryiGuaBDCNiewfM+b4
yWVZl7V7c9ITGY4nYFFmtomGPCGUiPmhuW4jfdL91fY6bGeECSEuZpjl+Vlp27X1
i66QNKJRVx6KUyf2ZUOUGtH6d6aU8pYqCix3GGHEBl7RyufkV4l6mDGubmzENyvZ
p4J4cydY02x6mpK7McHraCAMG0ErOkeTnSBFUbCfpDwno3jsX+oiAbM0H6xOlfv5
hLws0yeAoMd8de/ctTBv/GY9NkpVctLmitF6bZb19CiTbDNAsUVBHgudHVqCDV+r
WSdnrB9zPPzIlbPE5qzZqFUWr+c/Eq4s3X8UQVNQUPbfmCFiuTdyiwAkjzR1c3ab
gXBoYtkv1V9BI0fbQ0wqPWU+p8NZqAg3ri4OgIcCT7yDtvR8AEjS/PW/5ThWmXhZ
iDUkyu4sfbjyMAwbpGOi/HEwaMLCJrnoCGmsw2bk/dAdFfPLkQC0v46mgwE7XpSM
mTIW09qum6moRYzqdpGHgfUNyTIikNLK0RZv2LreH20xK33qBbT6s1RO3Af/L/uN
jwNqFr+h4Rvz1H0+m/hjC4yZKHrxQm2UEpG81MDJWPDqZFEHzqlGZsu8sjg9TcuX
A6+XAXPaEdmuegPX9uHh4gk19Qf7gpv6ulh+3Vwz0s5INtkWVC2u3SWBbaPhzU50
N/hQt2xLBUZdMns3PhKZ5aI8MxrSdkWFZbMWcE+K91kHZDcU8emf3jLC+zXe5y0Y
SNFwzU3M6PIONgSfahUMlqZkBbgC6rJHHWzR/EjQYWyy+Ki+TQmBoOn4LW7pxtf7
fCGjfo4p6wP3NngAwvO2p2hBtRWwL4sz1FR7hxdPhWl03I4LnJxn7FwMoLxlTBfL
A363gpADN4Y5ublmv1gV/ibrqjQUmcFcZoaqo+vQhEA81AH+MzqoMd/65S9+2gq6
bngPADAetvCYcLoO79U+C4qkHAlsIrZsKe7v+dWtPrUM1xWmxo2WuT5L8jjSVrnW
2dZsro5qL0TghH01hwUuomQJmE3jeN86q5JkMY3intvfBk8L9A697yesEyiWqEHP
RKUXBvlr7aNm/TIvCBUMGDT91qmtFlQOf9ADME9P/AEUtJ2D+zmNBv+hwYJ5l9t+
QNBx0c2tyoBlzcbnmKc+U2ENhzgrbOBkRT28LxsPrZqMSa4J2DLEo7POT2Awjk+3
7zUwKUnzghSPJWs7fL7QgVjdZ8reROmdmazy6g23eljw77XiOP1eA7bASPy2zwUk
0b205aaF1d1acuWjsUiX6Jy55sGL+6mIDRkTRdBWso3+K+LtZdlCmEPfGggL1QYu
hgyeLmXmxnPwVMdAgKHKBlyb00ilqPBhpEwqlDx1LO1fc+AcTcKkYWsk11lzKcff
EarXR2qAfQwcBwYVO43tNuEsB7FyW0k91P8em6IvdFXtlRe26ucYb2eqsFTYjigu
p/1g2RewypzWd+nGTYmK5nNb+2kM6DSq8a25xK3bJglhsOWWgi0bsLEq8ZE6zZrk
FJTaJ/Hv9A3FrpoY8GsBIqOZp3a4Qe55029QoxkjaU64IFitEVk8VsO66LD+L7IQ
4GjgD3bbkaKp9cPQH2etKfrKfrwK+DNBmmjPW+FWVcVl+2KfO/jZKopUFa8ZcS5c
kP/lbyISCFX79l2TwSmqLkpkXWqNNbT6QpayCA9oy1QaZrhLkk0/HHs3sPAhF5Et
0ncEeZkMiIaP5JpUh0e8nwCF5M3ui2k2XwutQS/8mETgOU/DFcmrtx+MzEBXT6FM
hVO0tCsCt7hI/P0lKVShCKWqbjoYS/JVKXEkY3zdovNcAEOGByN5J35ejCK6Ej4C
quwxXgEheWZlNZtRrlEW/nDxCVlHAi/ojxzKOecICCtpJ1o61Cvj4EzVZXwMkGlB
mI5uxeLe2AeAjv7uK2HZ3kqfUBYk6SgbmxzbQAW1UMtTe80TamaUQSIzXcznDS1F
qgD2gAER+cVeKIVSG1jyBaeq9GNjsUI3L7KBBPxIQCJZ9psUEi5hj5pySikoJ9uq
b6RDUmjMk8LBvfS8irqVxsPBL/sV8tahmupjx6Vn1qpTGYuxtN750l5OxAM4KMu+
yuA8DOc9JrMfwg8v1OTPAi1g9K/7EfcEIoRJMuiI5uUKYO6yGRWUKCB0CqBGubZM
tHy8XeWZ72/T+Pf8ImyCQ5wk9Q4JkwJo2NKoc8qhKMp3NNC1EJ983GQplmPyIR0R
noVqD+2SMkp0oQYqheCMhKWQ/cjRpF1mPqn321iTpKFu77qA+qPr0pNOy3TlCCTg
mu7No+q1MHnLrxCnCT4EvxdijKunQb8EHQOil+DybGNYxH+zNppc8YXhkNR5jazH
dzxd3TnGnlnp9CC7uYATWLa/Ov4Pee9CkTLr91gRJqsEZi8jqHQTObV0rqdJMEmR
cnjUtyOAIVpzGe8TOZm6CRnTEYLQe+1aFfdtoe+bHlgyCM+36zgHbrLf1ES7Cqel
CKqmq9ZHAQ7BxqBC3AXaGua5Aq/otBPtnOVCj2CrlhJQdEhNzNrgivuLo5sEy4U4
VQX4QFqfw8PPVtg+8NRJ6m9FvYKOGWoAoWmB+8ggih2TxdjhQWP7vjMIjZ/6duDj
LF9aldOVNhxKM2pXq49w8/QvA/rCEgnNdrIRpeSkFJX0BWe/swt4iElBVA8YBmih
/FyY9IB+2BF4b4mx0ILwjDWBVd7CEpEFhzgwa63zXv+ebPgvG2B4c8ktBmPiQ303
2udeNWBpHyZk1qpZfkAXy6IjMmLWn2DrNK0o1mA5zFBJgZYkUOaEVEmriD/9YcSJ
9k1CyjG+58yYEPLX/FXQUUtsyCsA0zXnGAEbVomrigcqMDXnhDourUr8wR+I/kQW
bs96GgY4To0Wtfhyq7R5Gnx5j68Y2uMPn9ptsctzsE70FVjuF4XirNICVTq6N7Og
VYsG8A2J3rlp1K1V6NKC4EhUqz/mI7ygbJgZkedKXU9Edq7o+4/OMtMKLJAKPY7x
EFnpOJH7t8DdXn7EoGlJ6NGYGaNglDBNWCB5EzjUWYZf4oqhxxPAUUdiRIzuIuzD
X5+oWqOUXDndaO0cZ+R/MqH+L+wbK2kNnEVha57h1wbrA7OJMzh5Vo/YPoEUf+51
z2emdxB8ZPq6IfJZgAvR4Fh0Uj3sqdfe0cOXiDR03GesLCM7S8Du31YG+VxnrHoJ
gsx5ppOcd0GSBs7Q4YbtM18zR1EjcRub3zOC+TJnUq2eXZSqhp/ZHnGn55dS8mVB
qLQ1k04qj2JfZDqtqq2DzTMGAuQ8/htm4P/W5Mh3YAGGwoMw7bZDAcuoFE6+31xL
hsjgxmJPgNL2p/gepIGECIpjc4Lya7PV5d0UElKsHKjYh5X6YPUlsAEa3yDAVyWK
9dINDaWDXwmZVGsWecDlob06t7c8BzU4g9uO5YDcHaiw9oONvvhfYa3MRkK1jLFw
loGKeVEwpJzvl3oPU+CuTZHb2pLFO837VjEzKNhlm95Bkr+5YaGUU//I7CxzwAh/
nLOLWIT/MSIB+uzqIta1U8v4cF0O6BUxdzgADkxoAJ9UHbOOKRp8/iuAGOOfykmY
ghjh1b67EkE+z2VcEikQn87f0SLjY7/fOBpdz6DQgDgZ5VOzQYUxts5BdVctJGb4
aXNnzgP7a1sexvgu4AlXX1upFzaDX1L4iL0msOFtGslhpXwe0SQNjjnQdMxyJYmK
2Ith3/ZtOIzIijUO+xCSR37M+7VflAUacYbtzTpaHpEbMprWqD7NXCwIbYZLzIA+
pw0rzOMwzry5BxOePSISIcbW/m8N/o8l3Y9FfgzzzDEBPwJ21HRU/jpEqoei+uOH
Ni74LnMv4r3go/4xrxFsu2jlLNwI3B0dnoGAQjocTUj7mkZfomfXrP+zcPNz5ZPV
wcwr+rUsT86f7g8YFLsXPhtjTVxLUxm4TQi5wrsorLe3e37nE61tXnaMPZHZKTe/
/30nredpoC2Wxr8iMCVhOhrih2KOgajYbwZCNkUD30IL5bKNEtwlKxYKoPFiKrea
07U1Mh9B0GlYifCXcgcbNPdBJj7cxScCEqVQekMT0JcTW1FAPshYCL7vL9XX/AbI
bs2lEIOgo2IPmbH1Dor5ysrxQKOBKgZvOAArq53lYbKjOb1veEC526AUFi14t048
VZHVhgRU2oJKrEnUMJDncsc4iXDeK1Vk2qyEk8W4nVB90Z+lbAZiKS75rwzlZ2lX
WP8nduYt3sHm8U9uKhrwbCKW7RmivysCgREKbVPcvRmdUc+4yCiTUcvVWXWpAaRm
bR58IwIQGsA6gwrjdqUSGtwrVfNftEfejOf5yLMWhkKDMh+Fk2cdrrFUHMCfjPvP
jvfS4+FZfVa1LTCh+Ng73d/UI4bQ2E2j5xh0OsgzjU6fwxZ5CmO6Hw6NiM5A2PIj
8g9aAtYnvrAFOqBWZkgyq0vIzFUZsg01K1IK74S/tEkqOVc/qgMNsvNAcnHQQnvy
WufnOO6MDK/jd4epxz6exkQFJFRWMmcTLF3pCogeVb3PJTtaBeyKd/o7Vrt1GIwg
B1MsRzn5VXdKLLSK5JyyOX+QwULbAAxDnEVKnPzuX7DCdOIz/eGFfqGNpx4jemsn
tr2O11cvOLoap2TcN3LbH8d2u2FO4xKnu7Sb0QQIepGHWa8rHep+r29sUQTj9ytH
cDob/3/1pxDZHFyzn7FmSu0mJ4wZZ/GaXaK/dwuXcDDQ+MceIrNrpD3KcmUIj6vf
7XU3D195AoebfRCr10Lo6KcW1Zd6plqqxIALsBTJWPt/RQIT3vtkN87Fw1yGRALA
V3nPFztyi1J2gXxwgKk1hT5KX/sVQoNmnOTlJ38dw+32BiLa8IspEVFpsqqesFuN
JXf5so9EsX9C25yu+wY7UemkHPULozc091LQ0aZc4m3Ny8FLAZaaPMhsy35GRxGe
AyFqsIFBjnfsRoGljx+RzNwOeXFZrn8kLMkn+tHHFq23an6L1lfPQKgqYfxnDu9l
vlMAd81jCoEEhny2SXWCwDDXt87T3kBuAKPXEeMzY+5mY9FJbAkZAwvEAZO8oI6B
hlsDIk13GJgjONEZ6eN6gJ2zt0h2RWNVK+YTcejMUAG9u1MNzS/e8UQL4mIkhlxG
d9Vvj4vo88RZDCVi3MTClFJOCJV4cpd3OGbZ3j6Viw+K5duovF+NLGQH1J3++prL
hEWc3/Wb62+hRmm/MUSioJ5+HWCkbIi+e0oflb+88QDdOT9Xioy0T2fFV/qkjaDH
iRW/If1M148hfisVBR2/AEd2qhpByENgDalzlJM58H5f2lkaCgUQVpoS1YWeV/+W
Euy/j9FSa+BbUyeXOtxY+qYLL+neUCijoKVlQixlGtjPujwtmWV8BI1JoOOWDjcN
2JmztjsB0Arm+wYojt5Py7rf+if5wl3rxSARQ9Icx6dCbvDMM3oIurEEWFcPYr8F
Q1aRtZzx969RMo6B1WfNOLg63PR9ZyGcjmpfdEWrD0imhkQZZSx0xBpM58dSGpQ7
kpCCAS+T0EqBPW2r7f/X8dKCsK/WqCRfKMf2xuNxf0aScZWfPXKOnLD7scjlGJ9w
cRY3LWOPnWp1m2DQmpuKp1pkTJ5EPUYVfI+Nml1zjN4R/rit31oZW4Ix6ZHdg4Pf
OXsU8LXrLaGrupQZAeCJ8MaOjSwwKeMC0Kqrwz0X7bDV18M9VpgVFnLxjuVMBXGl
o7wnj3RQgEF/qY+4J0HgeP1SuaL7IOO3Vq4cDQQsRV0wQ5lnyQqpgf5WfLS2LX5k
vUypzBSmA+ClGqgYU3VIfLuuzZGpucIJAxWPBfFaMn0flsOo+ipFm+4aZh+ulNg4
hn2xJHOs2zL/HG4BcnRPDbG4xNMVZbSuDbnLwjoRGjW+adle3mYNrPEWjxkEztVn
5VIXJKOI6e8ZFgzfrEh5p+fgWEErHq69bWbx4SI6+tVl1RBjRRsnFDM3xFIUUxx2
rO585OsqqKYz333XaiPbRuPJyNtmDvXs61EHLdThJUQ3/0sWGxr2g4MEEGtUpPs+
F50AzbpH63UtNlSvkXxpzTSah7AUrzovu+VSMrPz2G6b/5rTrFDVQEvYNTaAf8K6
5M2+eVvPyd0xv8jQ0Z0In31703OIQrnXSGu/vw0af6eHiL7y7jsoYXsBi6kvpv+6
NLCiqQNi1+HzwV54qu4TDiQSkarvIuINAlqGmcWVc3SukFm8NK+XLWQB+GkBLsvQ
pfvw/lLcHMyDGniMT1K4kodTDUtlAVqWx9BQdzzg0hmN6qE8VZOZdNHcR+yEO9r5
1QbDwieuG9QKzoiKbTI1s1TjdtwGbon685AB7f7eOMt48aGvTWvCiHekRHey2RIf
4ox29VJF+MJPfu/8o+RM7diB4QmAFXV58mztSkvGCDs5OEu5AbQ/fCZfn5fAOZe2
DnPf748XnpzEwLxIWNXPJXZERZxPNoOqfxss8wknal21EfbQPqySoLMvN/8301oO
w6X/ekDDHzWv/VF5oKxiyLtASXjPQm/rtv+6LFZvFd52fcwWuBTAKgLbpqiXoJQO
mMQU9mzJ0k+uiYsjsLGQ5LAUm3wuAJe3EkznqvbEiogTVB1QRyjh/tODWu7c5CzL
QYxkrzSvwyGyJlFiQV+Ax6kxmJoSdEjkoSEEBMKr8dMURqgGBq1cCyZYKUflnP86
xMlEBFfsegLp166y4DRzT5uzCjrazgwIb6jVlHJGGGUz+5XzYliVpEyqp2nyAyir
w4bhmLv/sTHztSpeHXqX3QuaK3Hu7yr7kGSfPnGxmRQd6HDsdCptxFzbL/MFEOdI
z8PDXWLmrIDBT827acuE2hUhmCA6WutXbknp9TScktLZGzd6FlepFYDohzciFEhk
DEJMwKljuTqqqpCH30w6yoY7lxP6OPSq2+ym4ZJi+fVSDNG5fkPZtRxV9iwK4zhc
ZbewBqYJiTAGtQV0tyBmO2HOFQatpnn7VilQC7xBxuoBm1bcECwAude8hch0t/P8
VWs2VmbVtnTnX72TeuCU94FiWZf6lqnWsxDCsHTR/gjLg2+KsjF9fboJDyws374H
NrSqIo7HhXaN8QRx8hZOueMT2CqEz1GvVGs8MszadfcFINiHBRq1VK7HPEz0sMZv
c9F6gRcOBmUNraGJc/nAOFxgZ0IXHFTt6gZRrbATUQEeEe1itm+HoKOO0PHYJkhA
t86ceMjtt3PtiWzTyMmpImVZ+kBGJzXgpE0eEfwiGk+UtGapbZzP/KZh3s+CTqu/
WNb9BXplplHWkdsGd3tpqQhmFcicEUh+H+YMnhBog0lbcxEJIpUuxBe34mmJs4l7
4lZanjAZnutzj+KavoAO8++tqwLe/yjRy/uanH/RLiVnsw0lVyTWJ1bxBRlsvRJO
OAXkWui7nt5ol5EtEX4O5XaHDZq/lsCeD+NctQghguj37lj1UKCVPmk2wKvwULuW
D8cjJR/uZhGmffyOl3p6eAe6loZyDdrkEbqtTEqH5+KgTZGARq9znqMTHBOSkJaR
Jsck3z5copU2L+/+Kw2UXOz+43Doraw//K+dTGREpIOW4oiQ9z65gITX36HK54S3
FBXZZ/NZVJAoag3oEa/p3qF6ORMHJuVcBtI/mgmeP9cNFDSiHrTxOAdjOzL38lxv
VZUKJWlPGK77W38UQns4srp9Zqtzy9mr0vjcNkXlE7edA2HXA4oPWJmVFYPhn/pd
ftAUqJOGNI+TLeRXeQ7ObeSKkxoEE4aQ2bFqWpq+vqSYbY1U7hGFteE6p5wS6IgP
h0pqltGZxY8e7xtASZh57BRoUVjfufdZLZVk2vFHOwQVxG881B20MG/QEXa3r+xP
kfmgXi4CB9p2fa3NNJi5z/WHyuYOjwLqCh/a5O1b5wRk9vJ3SbL+UWSHf2Cb3NFq
6az5AooyS+/7ywkNh37FWbcInofzj45vuSWUK2YFKzqRAu5f93f8J1b727ohrdnj
J2elykOCKBzEqA22p2kyCLO2aYlohVTIFJevzqMqUxb6bsEOPpzRXZl/FSCnfMF3
BvIjAl83eHIxnOrmhFOGUNwZ6UDS2ck5zwWzE/qzHj5/ARP/KIz9KG6NRq0RTjJt
xJb0S+5xcUDboe9tqw90M6w5iVKBb6qCsPxXiSUH8hEtA5uukfxz1nPTpe4tEpxZ
vVsrpPZYoEYulBfwr0JNDYFEdaENxSPPz6iR/+U4hhQpduTMaCUy2GsMthES67GU
b41W3dXN52ASxwgdmzymFnEXHEr7r7GTCnh0PBm9CI/gllXz6V/8pxQ+Ar+VsG12
ZqCZYgRG4U9PDXbdHVANkPVci0OJIlw///z2Isg3EaEa84884ZnPrdzY1vnEFq6d
/ATymxoULtW34hYiA8lwoY8cs7GcuReUjMlXBD87Ma2MLptbV+XZ3pUNOhdfkn/k
zStJ32UXX+cmcBdBW5YumVb+GMGiXykf3eHqIB5m7wNIO+BUFn1A0L7wtduUttxX
T+S8x75EGdsMKG08bdD2qTKfK2CkPw62+WYC9iCbfrjLbmBsjTVwaVMFZkGgIEIu
cuQ5nTKQh4IR9DTOt6Q8rNStwHOx0HNi6O7JHsUHTupwAXKfaQNrCP8xi1sPmvTE
W/ni9YA1AcicSa3d7UIhsQx3xddp1gLc67mB4AkfZ34FCmSIUvFev1NM08wOVT3O
gxZhwwVXHTH5hD3h1uh/wsWpX1kLGXDbTdF5VZUqs+1/eqiWAettafQea9x+nDeQ
of6qEJv00PuQMvR/YCxyozi/2Hfz5qFE2noffk9ETf4VGIrOUlrjgEldrTz8wqqu
Qm5zleBBDIiYN09OXqFvLugwoQ7eGlPtRZsunQXboTL+k8skV8wCGMy0chbE5PzM
f5uUqwuH/w1VtzZ8bck830QI/ZWDa/lBasGRxjRnHIcYkH213/BWU7oaiAUrXcFG
iW/ACmx/4phY3FnGeohK4+Y/W5VzRvf9lSZUmLN+YD4AoqhLjda9DozTyNz2uCxV
ODUkZIyHD0E99HnP+PW2N6UmM0RfiE8v6GMNFHsVwYmPwVSedYh9L3EA2yjWN1Fb
NiSFXEw6WE8G+JVwjbqVmcGFVDkERPzXYn39LcBysfgqIs7vsplFPK6iqGf/fQbQ
cQToucQ3FAwLYHtc1oezT84keS3bhXun482oN9AoEyU0UoQ044/q6tFwx+iYZRS+
jmX0eO/khQ4fD/UUcQ7B5SStefeK1fW5Js8fw0DdT7uLOFwHHK6CxOcLy/yLW6h+
vsRqFDsAW67nt5a/LiIuR1ACvTndtDY/JWxB3crhCBwobvLa5k8omyvlrLXGznD6
gf9KGHi3qYHnI/l7S6TaDH0ZBvXZiUyeqhDgZYjWOIQo6lhj5pSmKZsgRRVXHTPA
ywhx6J0cIbk81sUpT7JrNgPgbWPMTcpA4CzdUntzs1dqsd2PjjeuVOr9WfhSHSNY
4p58TMAUqaMYsHDvnCwNpP7VRxamHDyJ6pROHgnUGw1cRG/ReoeVJdum09AvgHpX
hDe/3De/ERFUakkZyOdUDc/MeeR4PnFHCMWYHaVBfRDIhsbTPhEeAMvGVTKyLGcw
taEka+fJRTTneYbHwA9wsn7/g8LbVNlKow1IjJRLxFx9KOoTVcb+V3GVX3Hw7NZh
wuenCYPM9JQl+Rtyb93UEaJk147bQzYC9IAayGwz/9Xdn1WfiOIyKmZCwsaWaj8j
XQD2UvmPFttiQCWJDI0PxIpdvVjmz0lt84JcVztyLJjQJ+iRkavalfI0meMPEXlx
s/nhF+TTx4yOFrVsUPveDYjYUO7L9Szt3B1osL/HCGhpZODEVLh5HKtBLFXTe3Er
NKs9f5bD3Q/VbvhscE2J5TxKwRTGC31ODJihdN5a4WB0pq1fx58utDgbxT+uupNe
vLiGwVZdMufCCTO1aiYrU0So8ABvBwBpaiI5hO4bQDZtX6uYSx3PLLfFVm6wr1/k
oKQKUxf6j0y96m+CX1LwQFQHIc+t2ZwmKTKmBXEhIIon3TE3hUlhYazIrcrfB5nc
8avnWMOaB0C6xlQO7wkYQGaXCOBAATAZXvkydlteolM1zEw70DDwWgEqtp1rJWxC
qTzk8Q78RPu6MnVAaAxbt7v02tsuWxpY50yJ1HxnVSCIUWqwRlEiWzMPbZeRYNmO
6V80wD5H4mq5YXOxd7jLgjFFlWtRGcZnM6+srwLLYmw7uGD/ylj0gf9P7Vc+EnYF
bca7211np0ZNzVPehAxD7mx6MvgYSkLHxnlOuFQw/sPdQBX+FpsTWAEuHsoRsDmK
5KXRYLZIuK6G/B+Tc6uH8DQldSrmR13x/Uqvyl46vz9BA9x7bDUyDyNGTAjygEYx
9K1h/RAR4k53BPhDWXryxM7leD3HO0P54gdetN2QTYZxWbA3+VNcgP3c+l1pjNur
wk5A+//tnIkWdC8IqOKuTohSMTtHtU6aQZ7vuVQSGxJfjp4KhfZnYzmejsbf5wPi
AhVFC4I8SODjhEuOf04wJtmiijQ+QMSSWvHgVfoG9aYRray9KaGmVRhL24YgwT6K
GLmA9Vr8zE5OELBtNbncXmUMJB4QQugNB7xqMp3EHQF56fksQRtO0f1zo00vhe2m
qUV/8KBPNcfuf41EHP2aIqPh0Etw12YeEOyaivly9YOa+bHQoZjDCozf2KghG7SR
/3DeaUINYIJSKWKXpaMRimiJWY61SswcTzfzEBCx4UvuqyjQdKgZ4rBfOgmQPbZ7
npbbaM3p7ZrQTnlTEgUW+z4TFfFdpfOjixAvNLH7S02dBlyRJOnhqjF7DZ+sZB8E
PLaczIK1ciz2e1WleeJorkXKq5+wYlhIGta5+uT485gjYl+Y8JA86D9nZxTeVsws
sybd6X45bQJoQTAIsmZEIXaQg2PyqZr6RIGEbxotpWYnZ2yaQgDa4Orlqellyv8Q
SHn1NvjCxVlwfsApeayP2otPatIHU0hPyZUA6rCA7goKC7e77yHBSd8Gs0wBTIGf
Js9W5fZKRCNeSKb+/GkymRy5nn+9MJh5nS9qos5/jltwTs4JCu4tH5qbMJS0xV3c
y/ep4sA/KCrJBiZTvmBVt1TFe+hpoDdwzeEh6DAOHZoE40c/IHb1NI9I/uzrJ08o
OVAAvIqZl+UAcg6DHRkPI/ZOZcbNdtJrpZloDLB0lhieZD4M6VGIkw519h8ap8GI
sbGa70rFj1U9F1alX0Wgnqfw9n5+X7qm7EpEADnmN00AAh0S0xcvYYgYFtnVWlZj
IjeReIHit7UEbwtpANjuwYSuAxWyU6dpzijEXa9PHd0NykxtKpOd4u2bj8TbwewE
63l1RLsNDHIZLEGAy8J+eJfVOLDB6IgKw0MkmGVnoxfVUSsJyUXDACTTlNSxfPuk
jmZal/q732KvAOjZHJ9wAoZqMC/9YgK2la0nMERmxMQDBVmpeD5qVkSvV0fMklv6
yf/HgbWMMXaPAfUNs+N2txx/U0V6ZmPa6O3YG+2cCN0MTOYZHUY3d0cPz8SGffVX
SuK6R8Nh+khdcRF1ZpIUcVMTeXanylbQ7aWnilWrrgPamQPCF21FrBiSYH0PxsSS
/7Knx2UThzxnea3RMdJceOWfhsKisyTV9bBZ96VDRDoPiZ0JX+peBqnkTxkzsusW
irdwiTjIBM2bvPwSsCTeUyRki4mbiaVN6hEjmI5QRCpYkjxPgt4HNZdEO9sWGX3+
OzY34EKLpsvfZwO3AxyUgWh8d499BznEnZH44lddKlXkBzb14RzW9QvUZToj8uV6
qd4OghL3KoaPkN3maBAQQS4tsTD8Q7tH1ITQYNZwGVxU/ZErWXvBu7uYDC5bhT7J
+4tDE88868vRWa+rReLeb+UsqTvWz1dTl7b5zR93NteLmqiAO8tgIG+Ybq0nxUVl
ywh6laIsO5Gn1bxvlv7C7AB3xVvrnrpYsASEsXrovfE94+eGlm0awem9t1ksBTZ/
/LC8q2zq8lgDrlXoB2avxGtKBLqCWHGmR6c5ErepQNegxCiTE7ADgIEO+zCMLeKq
+/XOLn5JTC8wPAhVEf2HFz+TJZKOz2E9ygn/cR14fdvdQY0/R1y3izmZxM4AoBvZ
blpj0at+bMxRllhm+mQ/FIqpoA5LwotFcFU37PpAM83R++FMX0MU7mDJTbR/HPg3
ThC8fAKGp1STIYnjXwZ8Y9NsJFIgrfI0XPfVycRLjT3bH+wTBWCzT7Mwl16mx0qY
V8HGcnvJuxXiqizXz1ooZgd9BdCdpyxOPl5NnvLbNatBY2V04MIcgUibZisRDIOD
vMqBrFT+1I0P7+JkUjTYaH8PdiutyzOC760aZT22/aT1mfWQFx5zOcy6ZCEEJ5JY
7FxQMBsgq7vwXSTbcqa4O5WK+ZJsditv0V+rkx9+iJ9QjjyBn6fqt5razqUUIMag
a/+f0IiPkSXHx7eD6btPaCmgOwIhyUckfCuK/RkJyGHYEEEFemXtgiSwuwxYKRKL
9nyzHl9ui0OgUNm4Ar4Naxo49+tRJx5/roarQsKqwn2QVZ8jZ0WXD1JqP+3A8erx
yItY/4XhQrcnr0CRVPEpxZ2YcF7VI+aRRHGxuKzVFgTKJk8vGB8awrUQqdUe5Hxh
gz+zHddeVvNI6LxToCG7f4ZNqI0XOSIdWRvjbP9r+q5ZfRnR3Mlb78Oj0rGpeA/q
hhvnpWOlRQVSdeyqxHawMHDzWC5kCXr4CX8zXCw7FktZYwAIgZ8yzqjV18PY8VQI
iPg4VA6pS7tT0iBowos/pVygMuZY5Lxads10njohMtUow63GOk4ba40Qff6Z4wSj
mGtmAHva0umuN+mRhfBRCouSvAIRKa+UxQ2+KMMhpx0auDMSKV5UUebopSCmykk+
h5QaOuOUV2fdJzrDiOD8xcclZwEOBYZyjSxljVBtnstEEWp4jDvo/obmx56IJqJ4
otHfkRepURUPQT+STPRKK7lOoTfV9ye1IK+qpKPKvX56uKmeqws3Ucb5ILiurMEX
zdm9TRubFXspqs9bPUgrQaLb0uf0peQz8Gftd5MZsKY8xMIC6Pv32IJVAuNRFdfQ
bdy/q3jtAxXYpBYKuSeglOKESMLq9jAPPytyaxQpDu9Dq0TZzhpuXktjxSjIE8Pm
R7u3FemVQhme2S8dFQCzNO1NvPfikZ6/rjDIkQa23MIqQuFEu6A1gUYjAITG7e6j
2/2gxXqn6T3h70v060Xj/RxIin08Yg5jHeECeZYiizso2NX0/YTlDvzd5G5VbE7r
Xkdws5gpVnA+6kAXfqo6J7t/9hQwLUl+0xd03DDqyv3kn3mAdCv10DKAVIXYtV7d
RD8OxwZ6nV0yhOv7ch+pv3tYmCB2p2wt2M4FwIrjdwi9zht9u3OpoQ4lVZLrJD3A
2NQh7tw4PkfSJO5yc8WOyLhoPlTw09UNfkC4+Lsi4P+rLLeAqSIFsv5UGgTapmEq
bvl+Ka0Uv6UA1v5oxU7hI8juWSxYGXX2K0yHskGI6/4hV5Y3mCN1i2b5KK3ZXTcv
rGOeb2XQ1N0SgtHI4QO7Zg5uNkABZUi8dPeZmpc6OxJo9LjrpxDM6oMXIPmb0c9t
PM6qTMm15Q37ggc1X+FjUIdpZwDuUpnn5GBXow5D95MWH86MU3Zc05UteqKbVgvA
IUJ04lbY+fA2tDQkuAgesDF6JS8tSyHt4ELf6lf+GBB7NZE3VotUnTCL/Z6ZBauS
BFNwegBbaIDr/qeX3b4+SR53C3BNjGgUf+IBN5Axx+WYruHV4DPfXoO84z5hnxth
upS6leGkQ84BsG+Db1NgzSrIBGjqroISUHI+OdvU7XqpFSt674ojyJRecyEp8e9p
pDGjIAFTW0L6aZVNY7D7yWvyef3er6cTw1YOR/AK52Ett3l4ias3tNLDewpFy/Ss
iylk8tDqml66RzpdlV33c764SgUk2CuBXCvedfKtG43hdYeLL69UytBuu4liAmIG
rINKJP5H0zBEUzj/AdVrSkUQA4apqZbOz3ehnNkWkXX0fep+9jsc/E4Vnu9ZCqV3
EDfeSwpJsO3CfPeBiaILyP9av1L4Rkl2JC+ViIEbP6Bj75Z5k7btX6hJGc5UF1LC
7RxE9XcpOsM8B6tdqVKDlAJavC7RYSlomYBcAuoBMBS6h0CkxOsvu6+UCjDbeA03
Kfy0bhxdQ3/CmjjelN2jTsGukJ8xQd95lXXi+CvRgdFnwNjq/hmdFDHPF6ebusG5
XxqGvvX0hBYyuKXjX8zugKtVEW1n3J88/jzsvPMiocFvpNVcODoDdOAFlbZpvBH1
t+KQ0mhrS+cECkSinuANCvRny7EWlaJ18NQc5NRdNzl5oVjnbx4CqE0YJ5XB2vhe
V1g1A5MhVnSYwrAmovojt7L1mjyv/umcpXCqojKEHJgOQStTM5IaScZTMqaRqfaI
FDinN5xUWomeG+lQm9tw9Gempn2LllchEX9XAvDq4aHVeG1sFUZQG1MRunrIRyEy
NcWSv9kwiM/dzUn66hIhHWeVY0wHw8g28YTA5vMBBwmBD8FLrA0CiFoV1Y8iEX2D
QYsV3edrQCPqUd65aKzJHYUqaEinYSUHaOQq6CZH03e51Txv4JaGBjbgDzfhC5t2
G45zU+iMPRMfEzTtdxhnlxVxeT2c4Osss7KoFJ+aNUC14U+MY1OhMoMup5AI5s9p
uJ+ufEsJhPRNx3gFDZyqG74AcQI//mvoaT/5Cna3l2qcuoE8L6kJYXmeW/4ht+tl
+LhBMkck+Scehcn+8YlfWHuAlb5LDBss7RCWo/fUMOjoYTOOTF4RascRgSS1fH2Y
r/W+Uvk7RDuIlDEpC0o+Aoir8lPXeGRAjQiEDzzrEF8xemf9X9j0TDttUXm4twD/
2pJUsHGle4IOf1bcW28UnO+8pMSaoHSqoVws5EvP0eJ4fzOczOqGVaX+vZ4jqdNd
XsbLDESfonG1+my8UhTLhH/pzhwmMd7TfERrT6TuiTkeEaulKiVS+8taDJLIBjbJ
D6BNt2x8xnodD4CJ11BBxdf+P36yXX7gSU3jNOs7zLByC36t4ldv3fDf6A4xlgn+
691RPhzzDw8HV1NmuMQCjya5hFgpb2T7LfcIq2NXOmyjuw162uDQB1AttadIWUwP
9Eifv8OrZe5CzrwhMbURMgrXNC3YPCIax0QvAUdo2294KOX/1UcowWqjMJIred+I
xiorPrWO327iXBH83h7a7QLJpIxvbf24bKv7gr0c1yVKIrmMpTSdH8uWXkCkt9Cv
tIhh1uS79CmXxhbYzaPfH7f8hNualbGoC8OzUBZgvCFHF+Jq2LdI5hpQHTnDgXMd
r+5y/f5hYdGaxdtlFyRlswNpF1S4rDE0oREHd1kdM7eh8iNeb/lrvRNlp9jPGahu
eWV+LxndClaDYvfTxyporQS98PKT4KQOX0yINkl1f70QqqFm7qnTjC38gP8pX2Vp
UcTE0lcWzJmrk9eVphMqW4RGNygGUiXAfqx6azw8BEmFxKuzVkGmvSEvGA8HAwVj
vB/02lJ5EBRL/F33+W7IvuMml98CMn4vkNIPEvTEbj131T0EhZAatPtAuygaphiE
vIyfxPykm6x5uePtv8XOLbV6uz02mKU+RByh9EjK8HTCXmljkod0Zzah74q3AC1b
xGQiDq1K+fIrz2M3Vp4FfWNg9h63Q8a7KmFiraFoDOLtTW1kjnSZMGmAxlgPtvW3
WRnkrj+rH1xKJ7TNFkbF2C5m6X7dntair3/xVMsY9h9D5DSO5mBa5b+1WFK5LMxV
EErLspVlj3dIddUyckVinHxqiM4pk4oe3E4BCuAZzlEaI8C4dzCQ5kOsmM2GqDRO
h15m+Sh5IKzp3Xn3W1+Z3lDwXwNhzrwu9MON6ra90KDAfkUYd4sTdFXG006D8rcr
tLlaWnaCWS5S9ELn+dOzfySh3+11UlABKNlotypsZQ7MrdPOypCqW1WZd+3k6PVR
zCLjbZKldR+DHRmHqIkL6qzBgTQHiQMJ10JxPpuoHBFqPy/x0Ndm+++O3OUwo9fl
PfgChMdBeLzg8LE2o/lHeEo4xTsG2RxcuBqnQ+NnmnOsughrzym97wm9sTTN9h/6
ZUYU3Ti5nqilPY9oVUQa75c/OlkHf3aOtWGcpVCs3PcvPe2vKr6MLd8H6POfoZDi
pm2jzsgu9FlOyZA6OeD14zCNQ/A5+3+O+4PIGaHgPXBSU6RbBeVuYIO9AXCYS/HK
USeMT+nhdwUtvg8jIm42Qydu09Yec4dt7S+SEsspML/YH/LjgRnpDL66qDUUVQ1a
Sfm2mEAG370SUNbFxoldwkUTrpNkaQWKNHH8fbYLuhTOYtyXKoe026VaQABRukOg
gCkFNsbbS8SJz0ikXMijxvqPK6nZa6EtGo/LmpbBCkn1+RTzq4K6Sd9QsputBZg5
di7RQN2BN6lcs/gC84mhJalD/3RtFk//uqJhTRT6vfh9Q8NdeewR6+de9YwI0wPG
7yvb7BfB0E7BbSFLbI/oEp/RawoK12fXi0GKIODLWvFRazBsZ8WXfjDlEWAK1i9W
/K0lfugyDi8zcz0mKT7Wy47QrxQAvjh5k5Qk7u2DctBJeuCw5uVhYvz8IhQlCzyG
SgBI9ky/lPtyKjlpD1cM6CUsKupXLkShWHkN0hJmC5yPZS26rnQayj1od7OfAQks
zQ4UbpgI6f3QZzm6Qpm7rjPpFtpx0lA855ZAD1hMhL25Uro5jz9SpS2yM1zGyU0W
NHpuXSro97V/sRVfa/IHM5ZfmLfPp7IMfi7n/6MTbicp6YIGLoCLbmSVsr6la3Bd
7U8HPdFyw6D8BvbjoSZY8fZCuExq9hQ208le/U/V0wgOXYZgcW/4YHGVKGcsNglf
NvSNJPN+oT7YhuiTincsNmIMyP4gexiiIsOdx4oz5tzAAkxEmJRhDsracxTBMFFB
kKAvLU1ioD4qBf6ZmlKuB4yl4eA4rjPVoZAJ3YBnL+aPQnRbKIv9mVLFb59NaV3N
HVR8t/PLsX8xoFYKqby1c0ove5QMRrAF1uaL0WpOixRcUI9O3XA8/tTzxObTWZKK
HPCka+2+29QPcoX2lH6yNUVzqM2XWW4VactPmEdVd8ERY5ERl/89zzCC3Nfhq/F0
2X3Gt65d07kIAysuKr/OWz0XM8hTvxlyi4U0h8m0fbIhk3g+m1eq+GsCd9MRTsS3
ntxtHupVX5zDcL2zjb3NobcfgIoLBTDAz7brz2ZHcevvRIoExqNfb6kH19hmclTa
Fomt9ppmw8JQUHrY2AYV1OpGouYMduHfSEA6Tt9Zv5kquylU8xv2IOp/WHQqVZ86
gEhnqe9n/ObzbFuQDLtUDRMfVbM2rS4SNN+83ZyMNEopXO9LKbdKyWPB4Tq2NlBA
x2UXeE87vFmsJG5/xFiu+I8mEzh0B8UANJO8UUm7A+wJfXS8ZgE9qm4PGR/bA6T6
y/8BLyqjmh/+Ap//lDjYTTY+C/hCDhto/WVLjfakL5LNNjx/aeZ9/II7GN5OlKDX
F5YZJgxA8RHO/LDjk2O9GuGjFX2w4uBVwyzOE0Di+MB6Ky0Lw+W94bCO7KFKI90u
0X2MJ1U1t0j/pI4VbRFWZOxqT5A3RCHuCGUeYol8q5uit7QoprlJsc6hT9qiWTwg
R0h/M6wGZ79wpLcyp7LGl6hExhUEa2eN0dCOW1JuY57CmCDLTkFmM/RMd8S6YwSQ
Libd8V4e1dx144s+XRAD5OYrHmnraq1W+LdVWfUO0Qf4kBrGXaDbEVh3xlSVg1rs
+o80UqQScAvsNhswfSVEqNm/OLnrG0eaDGOdOcMtt8tBYhzWaGrYBd1Njkjfj2PF
agkwi1zKHllAmpOxoSp1HUdDOSum1ZhWJli+G152c6ixN/hSC/gOs5HzaChBUAf+
uMWs8I1Y0ciGkvr45Bmr/xcYK6xwr2ahjFaOihUISqlp4qm8Jyc4B+6XO6Qnx4Mh
eGkZnmheUyjmkxOZGWEFKR6e22ZbsQ2AroBYT0TgGucn+8FsykVYBYygSkK0KR3B
bqOAAPWrJS5z2l+aE9RPQdjb8fFAzVGoNNhFPRXIMnSRkdIuU+2xzJcS6D5GiqFV
kDWbKyKIG3ia1TKgqjyVuLflcp+9n6c4JGergv4g23lF6c6YYFhGk+QwV8hOrlDk
/USDa0swjGmrA5/vQVhMXUBTTN+lY4VVul/yT/SJGjvbbN2KEkwG4D7QUJqQ8tEI
KpZgKDM6nMSafQ9GDWWUgMQ8xHzZjQz69PCZImWXoANmJeLCsZtlaKZpJI1sCQsB
QeQsQfJaVeODdLmvw0pKh2D+IGuWoiKbfIZsjBk/nStZJPji3qiyGFfwYz775ewG
ZYBKQYKWPUsSJBtYbbxC/st49LrTz6qKyisnTjfHtCRysSvJuXWylrtmCEgwO0Mh
V3MUESucYrrvXt9ACMiNaJ01hXfcT0GdfjesIZxlPA1+cy0G9YZlSft4N0JWdU+1
Yb71w/6giyEq60Kr2s2u0MOkCJuK7t5UNEAeeZioz2uta/PkNL47sdTJTnyzv2lc
kxCoUCa5dqow1vQMwOSouREgs7N+RoAHatXVbcPYSou5RPsHqcP7X+C/M3YNC9mt
AX+jmvqIbS0sQf+7RRRZIPWScRUIjTkybkwAvM/H6qa4/hLnwJsY/GejUepp4cBN
z1U+PzoxwCITLNXlKYN75gJON8YNW1+mup5kqjf01LZCoGUyLCiq0kwEcE1s548J
1JPuY5eNvKrqe/P2EA5RZuiJnuv6zmhjcBS/KJ5xn+yPch9gIcq/voXm3fbzPvOS
idFE1x9B9AhWNKfyh5LXMGERK597PtifDOtgs4GwTHFaJCZ7M4LkzWdrHhPMOo9A
rXmdnVLOuPMm8nH82HRGJc5rIL97Hfh75QaL2xk7dQesPj7ZnTbeL078toKNmI1d
ulsEuD5ht7rELRDBBj3xvtaDdpgN2dXX4aCzICU/ZYOIEw7SejLls3VB3rcztCGj
M7nUuvPxFWskGBn0NklkiPPsfFLJWw49QB2E8paQHCRPTFs5/0+m1YkhiUaZ/B2A
rzl3LOoBox0PDW+CHon4iviW81DPJuAC6tiEWYdrAGGJgrMa4NpSjWS6+P4ku1Fv
yfQApamk8uGVY9Uk/QdJXzrD/si0aCWyIKB0G4XK9Un1JTzPZTpSevvP/fDGUTJq
nfCyHe2va9L8Yu9vl0uXp5/CAAMQIOjVAXr/cf+Z9JEOH0vjBBBze2crSyCfvPTz
r8UCD+1Ary9IxH6xgGCiYn4+Do9VrDulufEcpBiZjzB4o2xnbgFHMOKB93MIY7GW
iz/UyuD5uA1okQXAaE5XBYBuvF2bgAsjI46vzXc32EERt5W8D1JCYDYR+jKFTqoU
1vabNzM0C18N92M3luSiD1AZKbPhwQnJeqlo9oVAED22A3ZWmungKjQUnIocRSbR
nHvuwwpBTuvXNTRrNX7iMN/bJpN0hIYXTytNaE6iTEPscbSE1qt4nsdC/F72rcP2
ndcODGtBeQ2hS4nnYRrf5MC9lRVDLp0abVBr/jF0PwClSGDUxg1tM3lOKO1UxR/r
JVb44gZBa0bAeeWVYBlC+yQTNy9SzAcNOhpik2YV8gFQPbezoE2qDD0t7CQXKpG1
Fhua+l1UG/m57EliUj08b1vIdDm8veXvDwc/8mctlyI9uDqSYw1w/edVFI3eLcct
30W1+QadFOh7/hPblqpK/kbX/XT//50+CzQct01dCXO4Av2wA8+oa9dZ1FbIsCTE
rXsY/7KbVyv0UtLojpOzkuOMEVs+iQL7l+3q8rXMAV4kTlDhrZy455w1d+7/mDOf
IY5Wz2cKBPhR/PdAaLeNroM9izFnPAQZgtyNQVqBMqJIcHcwr9GwIpoQUI3Bujud
0RBa1hgJnL16EdoAOcsVS2I7npQSJ3HCVncWUrKqq52N6DmId5151C0xSqTBYs/v
sOV2xFG1iZodl2QaY2FHrKamGt1nJB9v4WJaHrJSFYStMQWj9GM7C+psut46VkC5
4lLJK3hO6R3iOzysj7xBTkbT71DX8ZyP1YrCoUAea7x+++fDN/dpNdoE3RccHqr7
8MlZsTMO3//rwWbkRJixkaA0arA4ujpBcDzXPRTfXEflyvokNuD5VBg4sDRWkgtf
6keR8O3ufK7mdStoTDiTCA3pt8hmL56pWll56e3jqWLFr9z46NvAVGWERdrS99eu
UyLP8xgSTXwYfjzr0upEK4z19UxtVM1357oJGOaJjhDlmzcr69jHaZwsewdtvyXq
Wg83632tHhj3kbwZ6uWyPOJMhA1QPCQEx7Zetgb8edRkjm2N+OK8cXYFY8Mn+QHT
8lmBqmYHujORlL5FXauMOSG9hrKljE84dFp37VuBEpIi74e1k7nMbIQAPqe+G79s
lmTsZA6JXZvwDQM+DyGWO9rqr5rU+tl6BI0jdHWN2za/xSfNPhVmKhtCKQlMU7qh
QEK809hY47gjM2ArfYCnNqSj19hoaFmVBuM0iyUP+G/lFeXps8CWlAVKqtKvsHj9
4RsTtYn6ITz7sIxiN0+wc6jlJmeLg+TMxA6daibroCF+c8temFPjcls71GBHvJgW
YROUVQYny/DVZvamXjhDne+HKSl1rykx3lnEYzcIuUmNNli0vRroPVe4hfhD1qE/
eveaC5UE9/AjvdSNOF07RRcj1LNr/gaC8BHEORIcUEZVOuBa27AH4Fh8kBiS60LC
LLdGe4Gsch675u9bmcKWFTLen1sIq3U1IgAeoBPYyFhSKgIXOnnj77ej+uasROH6
G8dAp94aPm6Y9L/CL/VXY6ii3V2NBYA3p3DruJ4T+tGFEVQQqTh+gJPMkpdwgViT
oP0QzBrH6yJiEL8o+E+arhFx7pysuJMTQXTHiOVuab0O5t7+p8fHIkuQXJIbNaof
VFIe834vFx5XTpd2/i59PmLpIDm8Jtn/i4Bp1KpS3e+fOKyqJbmMaxrsn2/NX4bQ
j4FOjOVH63N3hr/bdZpJ7odZI2JDEoSD0PCtPEjNYbCFQNjMz6XlgczD3vnPfjPG
EdVi4S/3OIuUL39OC5zCc5gS/tJ13AMQTEt3QGKb5vumEbXhxZwKrwhPcl0G+7Wd
6aIb1MCpNF1gnPhyqsKRlopbDQvp9kocIRWbSkJNFD/oYCi7u/Ztbc2k7UR/hgxT
oqhxcdR8iDeWeV1D7DwVJYqMaFHg97gZYjZaipoLQnJUAPRl0Km4aR+KI0nNAKqp
lqdeRHPtrHFGPkT/bSJLb2T0Xsw4wzG3DnxQaxvFJBHc1uOjGdBXS5oGz7e0887V
k34yuh31QBfFGdor3eJOVU0jFN7iahzG/bqUm9avQ6h2MKqlMw0CvtBmS4L7gzKP
rYgsrvW8zEFc+drBuWrZQVd/azhPlAuZijU6vJqdltEpizV1XCXT0P54IU+5tVne
sb5MVZwSJkqEnZsd/XDER0kh+kFGKHQyEy3F0o7S3YSk2VPmqKsCfBi9iE7Fyhfy
LlqBuxmsczLxIy8WHIrwcoyTRr5bEaxEOGsBPo+oilcbH/1fC5EUkjpin3COluef
VvUFyeufM1XktAbjQJnfpJJR0Nw1h2gW9gVUhExOwMikrVJsdRcB1TyDlQFKeKDM
2SfDfnKrqHz8mPeMjeSxz+HegNyCbNs5uuz+VSk+yU6yt8FKu/fErlgvmRI+KvZ5
L1Kb4Nlqft1hJ0frRPNrblmxa6ru4Crhu/ZgZlp5TIRy6kHp3fIc9MzG7SHB7lU4
SidpR27xZ9oTvaWc/MSe9vNS+biEvTwl+jFizq9C2W/ZL5/0/KkPcLWK0CIZGFNz
hzNGEz0AX6T48CfN/hi0PysriNV3chxrngYJ0fENR9K0OncFy4NqzTCnPvCNmX8m
Pq6gm+Jdr/Yrrtx98FGPAUlU/BsVn9+TIzbApqRFncdeh3rcZG+lhBKhKqUplv3Y
lbgoZEkZgbLMaqc61nNCAAB6VZsfH4i9Z23nDCDpICPQF9NQW6ekhYCsDvX6GsMG
+14tWF54+vlH2cyebgc4b5g0sEFW6U/JMGKQ9nRtPORzVW8FG8188WmDM7z2mAaw
VcsDuxaskX7JnZ1GeXgeQf0HGhLhNEwKoQvYtYQ3WScxIuIZNfG/pEHyAEA+LCO/
0dEhO0tMsheZmaaPutVpmUzQrNufqQsRn0rKkdmkQPGoVUL2IVI8IRcKN6sldjPG
JMZ5D5oyUwty1+bbzqgn/kCXVVAp+4yqCMkU4UzANPQ69XCRIow+MZzItJK5kz0Q
7qj+0pLLgbpkcgyyi+RXUVi8yUp+Jcemx9kl0xCwPsZe6rzC84iSiGk7JDWv+q35
MZ7HjltnknGRrVSzECp7fjI5nw5onYKLRXU8hHB9zWomJHwr56oUZ61+WSXN0xtu
/NGOgBtf4kDN1RRqajZ29S7vIu0Kb8+W7SKYZHSKhmLrmU5k2l9SF8Ovz7f4QpZg
WybiK14A9BTwrCdb4tfH4yOVQIlgFd8oY4EhYI7gKGPDsL4KB3pb/cyDlA+bZkr8
Szul6QUKfRjCwoeiF+Hz+cNaFTlVVkJzyx4q9wpmnE9+ZxmPOu4heWr4T+mO0zJ5
m/gWeuS0sVMyWCYJeHWLbw4gObuj0cSY4rYObWI5+y+CIxyhNYF9Ke03p56shFFL
jBbHfVdczK8MaUeWjuHjwwXWqFdo1MiCiCqSMqww4PNgPvohaLKN655ZrUYLaXog
kiy2Fw8ptPSFtvHj4R0gdft88gygmEZpsDVVNqgeTD3jVskNID5V+FmnWu0jylot
VfWVUrf3X1SaRZaLCqM3KdY/PQYf5R8I9oOaWDdvEk/coXzv32qE76fL9AdQkbyf
tTXlEP1npC7JKXhJLVB1zc6C0becwtCplMj4wAar+ibF9UEjJyKBODBYBxjUJ/lY
KETsR5EDara8PSLMxfDmXLg5CRdNU4qauChWpi8LdOWJsOQbmyH04U/YVWL9LIxe
WAko4VwrbCjbu+go9zUK7OzONiUc8zzs2CUmlUl3Zibc6K3lSf7SY6uYavWW3pkO
oVlf8glziC8fPdCtpNu7lq2hf1IzU7/IQr0E9UGpggXOCL0Mu30w4TO/bO/pZZT5
zrJszH9G2IV7TkwnDMBo81pS1G1J755TOjKCbgbRPknxHnoTUPZGJOxHdzdoxXP2
rQSdJY0vU+x+oz+JgjUndIyD6SzNuO0il9KKJGCs9mLT0EY1z/foEHnyLnBx7SD4
m2o9dpILM+WAZ+uCFX7KzTotBiKc01qGBfYzhjNeMf8+IIEw5HUAX503ts1qtJ05
cfv6a3G1mtxxxAtPB8sxvijjRii2y+p5QWFUqwv6mTH8K82R7f2Au2ITIcKoL6Kc
keQxQ16pZFg8L0x0vk6KBUVI5Zamo/T2CJuBF6jmQcBr8FcfJcSDq4owWS6UcgKs
B1qS7nrcvjw6/+w0rIvAewhu4uKg0BOj1DIUM9WatJ8UzZYEghPjgqO3faM58OCQ
4EcM/6Nf3Xh07gXYoFr9viGFLwfA2sl+/6ZXtwHpW4Td+Xiqjx/k1CQPpAgruTUZ
eEZE8dYLdXfoBUoqysVXrqfy3TsLBssMPoNYDwg1t47wb0M533tvn48rMlCIH9Ui
LSUtNUQjTNwyP3oUVm3yqlNoQN7TIZVUqM7zIHF2swiUmlpdE6VuFVT5YgnidZyE
bEFvG7mX6HPPdueJ2F4ZjEXz0ayxWcQ1TA5WN7Ay82toNDzvFe2Ggtq1B/WEB9Sv
/5tWzPZD2XqZ8NbZwTwZxid0QOoguypm9vkIPvqCq/7PgLj/G0wMqbzsnli8keLJ
y8/itbYlX2dQJl1j1z3yO17Z70kaXf4xAXBCgV8Kg2RC3sBfS9AIzRY13ZPNXcLo
wl4lTIgrbGZ9f5rSd5LcDCfNol++64WDOJkJhtJhQvCsD567Lj9DYAK7vNPDlLqa
KTSNc3hMRJLhZlrh62YSapCC32STXfCo4r2Ton0+2AUcKOkVa9I7Wd+rK5KlCgZu
uwbek5u0JaKmctU6KIMFXZnVl9jrzfW8TjnDXPAiHLVJkfpEMQV9LRwLdcz+oU+f
XP6GJUvy4U0x7Bz1sq+x9ojeQsERalHqbh/WE3F+23J6njnPkNUyUHD5SF83I1hq
3JCKdpBZStSGZ3W4yp6xoH2BBwc0jd9v2EwxEQjWifXYyZbU2uOuzaYWG2hx1Sub
XpdqpDlHFVogZ5VZ2M+nrojnUxLS1KnPPhuD5OYwi1iF1BXh6iL9kcMGVftVZBTN
1aRGpgkyWADNi6FfBVpSklz4B/fg1/Q2gp8HzsCJg32hhxlFyfHmxxXdxobYxHRs
8IjoMOUtW8hwnwmpHlYqo2JqOdEKaWvEDoSi6q5c/kOmKm4puGcauFvxdbIsmXre
mxPhML69MX9TsYCOCDfGStOex2zKGHEo7b13OwJ1HOQFxMGh8gld9FgIIXY2BgFw
0f2Ljufsw0dGwkxi5SNhCI5hhSrIPluUxGucQr+x4UW+9FW2mfEFjTcAMZ/UCSB9
D05k35xfNlHu0MXi68A+Cvqoxs0gmBqo04otTb8USXWS1srXG8EOIqo3l1fe2o31
U2RtNpFngDnZcO8a7RlDGFy/0GrdKUeIa9fnn3yVMzREfaurFt0wdmqgdTML88eP
+ZdAfArqMJ+Mw4tYHdd/X5TEf5cMXgaLbfM6w1LFPs+hfJaQuhmp2yHkztcfjiO8
vAo0EhawXSiZEEh3xAJkpPLJDgyH4siSy8fuOQrWnfMR/8dDQoA2nVYPBoRMwtHj
4HBbFm6SR09UhAS7IcDgNqMDkjVzUyLiEl0u7FABxLaRhTgH9JrjUVn2F0Sep5o+
9y9lGeCVW9f+qurX9U58Qrt69cH6almTVmFl8KkTV27ORwtErWqlQdqMcpOFlYYQ
391/e15kOtxHel1SP1cupGcxD3jl1rRvCYwu2igXfHClZCYQRpr5EWAKVQ4w0ZRf
w4ClGj8flA0Tc3WT8SGcB7bErl0oIW1fLVbDYkqBFH5Ki/y78Bk/SfZ1nLchXRP3
V/kS7yBosm/lGLhsT2iM5iLzxhQe5Soivrpte2GYttagDZ5BEiapUF45M1dEW5uR
MRC/Evxv37G+HHMdKNye2sM/lOjJNRn6W8fsOUUZ/yoXlDwnhIbDSMgxdO8UiK8I
djyWatqnwV9yex9QhL3MQTUqXUSoTryXalAr/rJ4B+rLuKfyeg0omXgrmqLm0UmO
ystfT/IJMACnyFMTe3jUWze80jJef2TlqhXx02/kx5A7/RZ7/TfrH44gRa56DVUf
ghAamxGO7USpjiV9sFc6dmBFjNbI+zbRFhN9MR/hEsODSPf+4avOJzoUdQB77SNR
uYJ/n1SRuVgOaeFJ0VmAxSki4K+v8tgDEa3CpHQuYNBSbZEI4lBzrmY3rfDr5QU0
hY5OH6OIHMpSO3oAT28S83/fTnl0tTdz7tWVoHT2pQ++cyb1SPmsopcMqtfdNcCF
ruFpAZctVyxoj4/G6ryRK/ysV3vyudNdLKyn/mOOo4Ek8X6mSGEJyp539TQcbZkB
x01jvx4DqyrmE7XqXcVIqSSmapvonkwwmUdXC+WKuHOLYmGbX4DlBgzNKZ0kn0CO
xAwdmtOs5sgb+eTl8OUyk3jaq6LHvh88aHMxA3xEk/u5dcm52VBoQzuNDQlSabh2
7E9wa8/BM1XMASbN6CMFZts6So97ajVpnqXd+PSZK/HzRjgwjq9eg1+QFQHdt7Xt
iAvZ8jH0UzxaEcXPWPJuzmT4jdrPJBBPE/GyKmphUJh/LEMW01MivF3FctDRjW74
97Y7y0p50AC4+6g6E+s6fdGXlUOUY4COI9vVkDWel15qsP8Jwgp4cLrITc5yivpP
cOqi+SPiKMRkA3iqrPtLWPjrr5Pp/kazU6dfLWhT1G8u+BiOII6dQNdQTBv/YvPX
GwBabdTgGjVUplxURQvFNK+Owa1UMfIfHh5ycSOo5oyOjy748V/AUP65hCvMqnwF
x4Btlb9aI8SG/TLhuNAMVj77/qrlN5HqQh+MvUUeqxgsbhovohq+rwkoNzub+VUE
JbeQuwrifEdWS/95E/TC7ERDnxmjjz160V0JeR71YsefsI3QrDlH/nr7uAMecOro
r7L2KAiQ9kw11BHl95qg0YdqvrLsg8O/Gx43tSQGm6poX1d/iyGu6uVV4aGP4LrX
fyyn+FKaTedHMTt5oqNC77GeGMGsJALNPanXcQpn5OUsIfMDiAt/Pq0fwnY0ZVlb
KDENSFYPlN0DYVVLJMWxelutiIAJ8ar2XCwrGAXULoE+igC06yJup2KoXog1dRvs
maThXgQrNxzguanQBMTRQtHgjX8OkI74sIp+/aJRIuxgjH674ts4yvbkBE3IEyyl
eKbuNt9nJsynZBdtAhv62IYkfj6wGZQwgQCB4K9uubik9UIyB88/0Hji1CigZS3L
+vaeYwy/3bgjcdvKUO4M3DF9sVuksFxfoll1+HNMhoeDmauAcHiAjzAXol3CtyfX
5azPtn7q8ZU1L3y6yINSA1dEQecW1x1nsrhFJC3CAQSQ+Li+kdnOaXE1/pCsETdj
pPUY/Vc2QFEnemXRL77Bq18IBw95Z250aFTtNedABBiNyY7lI5ClKUHUaTVSXeRm
MJ6msLLhmaktNxgNnNKHn+9HK3BBiY27eKztX6XljcI=
`pragma protect end_protected
