��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?��D��@.N��w$k��&0k׳���͚,:��I�oü{{1
Ե
�i��qQ1��F����0������j�Ys�A7�Q������܄��j���̀=R�-_�4c��-��D�b��� ������	�\͜��]��xE�q�Ws
���Џ�4��[�4�%+���N� ���say-4e|v�j	w@$ |�T��f�b��8�f[���U�(:�����ye���Ű9�![3�[/Tl��.��ML��V�q��K�މ��a��)�f����>���\U1D������9T��`9�a�� f�R�a�`8�Մxs�ȴ�dK�p���j;�a����v��p9�}1$�����
�����y�z�ߙ���!��Ӵ��D�X݅�
F��h`�D˙n0K�kC|Y"l�%H�z�����j(��*�$ҥ��Ҁ)gR-��4f1�P�_m�֖D�F��Ȥ�#�Q]�y���`��Z>*D$�K�f�,�J���H�	�_H��{!~�tH*��O�{?�&=�� -!��.�.{�&�i��~�!CH��""<iD�J�6�/�}z�9��m� �
 1�6!Tǚ��A"BP}�����'��y��Xt@7r(\^2�"��{��@n�1�M��{�1t;	IJi#�e���N/'@D�}���92ܱ@�k��`jP�7�5v��y�g=�?��q5k!$�v}�bG��}�
?���}L�J��mlB�e�ިb ��eS��v��[�U���gKRr�5�]��4yZ����|�/���b���{�]�c>N6�^�n��##68��2�s�1񜧞�z��E�X���D���'K3H����Ұr��	�£��ٟy�&�%�U������P���&Y�����QFl���=3��%�>t���"���|��P���`e4�ٶ�^�6��Sq�_�$��E6�Ђ:��+��Ғ3��h�=�O!	���� �*vz��(m�G}�5��˪xm��큥�l丐w,8��l��Sp���N�N;��u�5�h݁=.��Ns�P&�v��J���i+�<3�ӷnO�p��{��PIa��%��>�$U\��_�LM�CӸU˹ͽ�F�"�N�կY����5��-��=�@�U��.�ڝˢ	�y�Q�F�|�v�aI��(s��H�i@a��kb9;6�-0���GǄ|��3-,6. ��8|Z؂��y��������y�@H\�v���L�8l棫�>�%��i�^��ͤ�{#�cC��-Ƨ��}d�H)��+=�gA!�A��������Fc+�ƌ�I���b\�%��T�l3ŋT&�kDS�������`z~�_[}���>���6ePq1޴�J��¢8d�پ�X#S+��@W���r���G&��Y�Sv@�����饧�y���X�ͦ SZ	��p�J:���)h�)�/��0�	�~O"����m_�Ag1�S+�:��G+��D�	�%f��T@���e
$�5���~�f�c��˟"�]�B��|��� Y��(gSb�\Ik�0�8!��0t��a��~ܕ��z+����B8��_�!�M��C�}����w{D�t��t��$`ۅF#=N�:`ˆ3-)Ibk:��M;}��,��%!�VH=x
���ן�ԕ5�,NQ���n���	�^��]��2_a(!vv�*χ�ݓ3���s̖��d*IN���'sà������P�o178 ��FjF�welJP���,��f��#��a����&��W5�ẳU��]=O&49
|Y�d�҄��ޅA\De���! ��.�oq��+��ɛ�u�!7�d�Olb 8��k�!��<�=����{��?Mc�����4s<�-���޶�/�G���b��5A�UtV���-!�d�
A;B4��:W��	����#p��3N�����\�!J�I���Iz�8����f���}�g�?@,۞jV}jn�g��M�i���+@�O�Z&��wҧ=I4�(Ή��hI.,Y��[)�7vA*�f\�l��\X}taAgD$f-2��i���~@�#L�B��e�Ҫ�@�`�F���Έ2���{\7�Tv���	�U�gl��c����4yS�f�v*�?��yP��ځ���ǒ`��)B7��ORR����
|�]�5 ��<"����ӭ.cq��$c`D�������j:������$CW"&� ��c�P�x�[��(���#B����و��E+n�Ȝ�o�2���Z�g6�,���$'f�,�v�X�Lf �H$1��`�U��\�ߢ�I��P�b�8�*�߹��U���+*������&�K���a���\�#:�0X_��B�9�`i#��i
'�;nûYS$Z"�ڤ���h�-��v�D,p�����Mk�ô$��b*,�/?]/�*Ґ�U;f����̰�|�a�N����u4BM��4��0/�[���i����̔y�Qs�o�022;7�}ᵙ��|tȥm�:j6�"�#}��04���6�
���WwA:��td�^~���=֒ZVkͯ�V�(�����x�J��?D.�@T�~��\/1�!�P̔&��X,�b��Jpf`��2@`��І~�$��8����b���z	��K�z���Vu�y	�ω³8J��s��4
���[�i�X,���*������b�+W��{]ī��J0H��8��S�J�An�soᢱ|���( ���WJ���b����ah��ם��$��V�䬟o`,�����Q���)ϊy�Kr�L;�w������zk�(8��2��a������J�1�o�8��V�ok��S�x�k`�ZȦW$i�Z���u>�)���T\V��JW��R����;U8�4�D��b���
Y`��-~��[z�m�88�ˌ9����,����qŁ����"M�^����H�eXD�*�g�0��5���Ɯ&Z��*���>�s[C���i_���[��Y/<Y����F�.ЬuE=E�'��� Y�P!��:)t/-���IM�����[]�V>j���|�#�M��"�F?UP��QN~��}�`w}	��;��;v?�4�ѻ􀀶�J���������鬚RZ����{-M#��`��L'�D[�^r��W�`�<ٗ�M��TwY�V�lR�q/P��NS��<�,�y%(f�]��o%����xCj��B��8
7�A�)�:�� ���-�*�ʦ�@˓ԋy��誉��[���AC�8��,_0�M/|6�@y_��I��_N:o��3Q������9�*�'��MyR�qL�$�?��-jvw��-mI
�e<ۊ?�(,�x��"��Z�#ϕ˗l�|&u�R{J���^lĠ3H(��k5���OBO(-��|�:iZ>�V�it��ӂ|7/"��q�r:�����q����k����_��?(�:��>f��	yhuz�<=�-�ㆸ&RD#���R�k=��|_0]�4��B��'�mǟ�GK�ͯ1�@��?|t�3�JD���=�yy��Y%y�N�ʙU!����7M.ʾ�`������L���d�/׈4��y@
fx�R�v�f}H�Yp��{lhn�ϽZk�����:�dC��b���d���e�T胷�Ɵ�$��HD�w�8ĸ��}	��}��N�8�_��7�ޫ["�d�]ww�3�3,ZU��1�!RvI&��si���k��Bu��Q%�kV���<ku���L�
���M_#Ὢ�G���Z+�F��r��!�#k��Y&��$�hv �X$�L�P�c�|Q FQ?4����!�g�WҒ�N	n�Bm���z*}��$z.;f�ٻ�h5|1�
N�63��]�3d^�d��ݛ_�q�7a����w.;�۩5��%���5h�\����~9�"4n�`+�Ʈ�h� �����k�D�)XH4�qS�c*�i�;��	in�6f�&�V~��B����:=j������z�������@�X��!�3���"�]]8v-ICuXG[��PQ�|�T}Ͱl&�7�����Z �)� ������ݜYX�0����-U��kZ�=)#!�f�K�����*F�>|H�bɠ����c�B�.j�1#4�䉅����O%�%�<�� �q�E���l1�3��0;���*���|s�!�{��!^5���A<X�|/=�Ѱݝ�˶Z"���.�V�ک8p������}�!��ÊN�M�;�1��1��P����+����