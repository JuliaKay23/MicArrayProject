-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Uy6k6bhKnyhpvsZ+KmlXsXJhK4/r1NqPOG0mbL5ViRFxY5ugLD1YSU48auhpJbve4eLtbOge4EGN
pvaC0QhSBGrxlo6KanMEZsD5n7jLRKDEStMs/tKxtUhV0W/zhVHIPPC09MYg9JO76SWu5md0u957
Xj6C5mmdkEp9KjxVGL5AoMN0XdnYGXf6ozbphAE+h1eHeHnzwEISLlq+YuSDkc0C3x4rwgiFv7wa
G//GOeyssk7ZaBHgOfxMXjnEbWUk2mNeBjJ/E3MNRiCpUFWeObk3U1JzUn/5LoXH132FBkhO5oTq
A7+OKEBOjGjpIu+bEbcXhLpCMX9lose3THWnqQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7696)
`protect data_block
tNjYH8jYkA+7rE5yeUGlgQe5bT6qrmk9c816axOoO4Q2Dfg+OMRIbr7iRzk9/XiLIAcgPswmUfgJ
OKJvceETJefMazTJWvgvrxMt7j5vPYDEo/hPD9m7vAm0bAB4LKlmcpYQMe6O+5Y5FfrqODn7BDjk
jodRiY3rcZ54qJIYqNyTwCbwtyUYvAXIsJuA4WqZAbwnaonKfuYyaE5pTYsnbMWDqbzf6epcBXtq
VxIx6xM/eIYRig59ASk2YLo20BHsCkBt33WNKbWPZBCza96cu9ftD6F/SMctI3CYeOw0H17Pw4Ex
/CmoKfiUnKtJN6GvgNZ1weeDhnH4RtT9d/sSm6gUqjtEPfuY5I32G2wsCHA5JMECzyebDvw5Jx+7
4zp+OSCWupNiIdWqQ4FyxjqarJ2y5QDLVwbpgmf6h+S4PriyeOfB7zoRscyW9UHkaNXDEepOc/y9
wYaJ//qwOGBKibYcv7VYuK2/kZkaxeeGQ797zesV0WeeRTZLHom/EADD/lRm8z2B5k1qfI29FOEW
bQ9jThmh4koP0n9PPX8FgzKFXFF9Fp734J/yiIddM08NOU78AheHFEY4+Lp7YYIkq7ZJXJtKoQuQ
D6Mk0a4GGfHRBnIET7qe4v6SXONrzclGxq+Ij0RH01xcLUwaNXV2LOj3+Z80LHcpJp9NFKOGmoWB
iOorNRNa5a+DWcf8m2vuRugFmWxJKJZO9DNYJ2NU0GlOMfQHO/ddFK/d6TRP9MwcOql70oqBtKF6
5ZoWneeXjBcOvmWY7f4C/VOvn1M2fYvjex6I15YlxbCB8J6THsmIlM3OizOOKe6ICtxt510HyIsC
UYI9vdacjBk0qXXBIi/gYtwWQZJ92WiESe29YdBNp1cr+aX+8Px3jfWLyzuStN5pkWFay5x1bjnN
xotyDd88b/tiAvUsEI3UGHvpPJ7p0WfN/ll5/Sw8+2Vl2hjZ2THFOg0wX2QhQI83nlriN7sNkTiF
SFYGYPzlYTmkSzDTJkstNCbM8p8wR9obbUUw8ZeRw35VAj+c3uTGEVpfwD/nkle2sXboV9ms+Ija
u8LyU653oeTFFn3YE5zazU15qaTV9SAOcmDSIU5QRlLUL+SQ0Gg8JXUPGa1IS42y1kHMec47brW3
6uBj8z1ZS2ccL50WMrzaegKhLHVFxiqCD2DJbE9McGj4IX1CvmFKW4jKGoQqlPlNRC7Ait4Nv0za
dFVzn2/E41DKK+Ds9sH3AqG3Yy10jeuJ3PrKs2bMmngBp4SrgSDKuJhWbsK6oSqQx4pIOZIFUSh3
LPg4egfzQwvJ7mSZIdpLU4T48l1BYB65Nqplp1zJZwRhbc7gaY9kyoiacFdTQH4AiqBmbgMjGtqM
JTN2epBqZxkcOKdQhA4zLAtzNG8sDqXf9Ds/iEcC7Sgy/w+7uaLK1skpfX5Ff0nCtqjf9V3FVcmh
Ior9eZGNqsQP8Vh979fZMSLrm7ewnz1s1bK/M1wNjUWijufX72ZIup7Pn0DV/NZC+T3z7KBemHVP
jeTkAAUh2yRYJYsgNjl9KIPBDh1FE/FOarvpfE3EC0dM9BihPtKst2pPh5u7caiSuQ+4Q50/KRDO
o3S+t7Mymi7xGePYRIfzYTHJwCp0HIjScH4OeA+zHOZOoT054wAjhgrWUyultUq2sbawFS5/DdMP
qP3wvj8RHZERpWef2uMPHUXaHdXwhYIthHR1w4xhZ+220fP7i4aGEHoFCFLCKAT+vE5PynBpn+9f
gXDXccgTwkPKbORmC0DxYFpkid90Z28jVWgwFyPmfzuAOJFX+epLoOAE4J7pWBju1FJbSiWCYzWj
qmfEN2J6vhlj4OhfPXJrA+31Q2/HX8mwdrrxkP343D8ByRm/Z29wMduC+97Zaya+9jMLV8Hu0p9V
F0nsr4S01RDjkG6GOhkcQgg1G9M2WvS0jmuDb95UkQNbk5EV28+W4meyi0sPizCnLZVa2ZKSOs/H
+VhoMtxnHfIut4o3ElR4ymOPp9UlgJCiN4lz5kCQir/9gnUQY3aaQKneXfxcsHTox3BsY22aY3d5
jrEOCw15yZyyAfMtz0KTJG4wnM+hBwejFFJCvVe1SsgsjgWlzcsfsGUJmsvVS7Gl4CtbdMORcTkZ
voH8Krj7Q7gEazL6cPkElro+NHxyO1cgVtoTzN3Z9rN+0f/jwhRH1i8ey/S/kOmxqZCTxPEPpx7W
aKxf5m+pDAwQ+1xKFiP9Ez2Ay1N6wUUaIg0dsKEkgwihdLO9Y8ZNM3AzMhJxW/z9OAGFu8vgJ5jU
7p1oZ7VRIpwXrd5hYHmWFvaK+YO7oso/LqUtr6BgHhveU27hFpA7L6Q2J9YIQ+w9yEWbi57mHbeL
ZaVuKJxvGabV4SDMCxy2CVYa2+X40q3kmrOCtbbhHuO+kSq9tIoLXGzY/KbP1s5HG6iDZ5cetOmF
PExelZ+o5fgmJbqETu/4OE+wSJW7wlKzmvwqiWx54JcWuDiuasLVRm5NX9s5M4hVuHPZ4zZ3292/
Miovn7IU4NA0V2PrhNpXT/vnoQ3h45K4WAPzjWDUxQIqbIR1jnzLLTqui/jAJD/MI+31WYikx9bP
fj851qxGOG4VpheJ7jelVv4L+SCjldrcc2Wi3HFH0QsqCh/ceAPE5PDJmgPu0mMr00DiJobRt/GQ
2v1oPodIdGlr5y3y//e1IArm86obd/TfDP3R9nGPIHivd2dcLRguVT7SXY4j29tDKZx9WMTNASvw
fCG+ZDxAHtu2D4PGUrSA2BgLmHZ1ish/UHUr5M3XQY2zuMh2mhz2VNNQvACZ4MrY5DnaUHqVLjmP
puGGAwM8+TYFlq52j/mRhBXZcjNFA4StknF8vy3WV6up00ZvFu/SHQA/QkjNqR+hew8+fYox6Y/U
yI1MMxwhN1ypsJ1efsaNFmKr6kBNlr981WxK5vKGHvvEdo7uw3tDT9lfy0b1iff+ocwnedkCYamy
x9go+cuBtMXHhb9RRAG4mYW594sqhyQ2lpC8bgKHbeEtP1JKEazyIFrn2DoamNXaP4rju4dpjzmB
eFuesCKKKgLXTTXkLLsFRAmMSSpOYyyO60H+/F41uvapO/ujRX2tVElZUN9D4nzGtJ0MkmGbj4wz
gScBFPi8GF1DOnTqTWX+H/MWzdnMYKmQkcCyKZQ3HhjtU/X9JGCCPSdYwIO0re9cwkT0qvwa50Tq
3s3ejT2gz144zD7HzBYQFq+XYeeWm7+FOy6rfubZaVyba1RfY8TvOUI5kNGFQJcULCuF5kt11e5+
Qdog8pqWQst4cDOf1C+HGtUtlzPJBE7gPSfwcuBW/6/vM2LdpLNyXSEHBpwp19SnepOp2z/Sl6Qf
r06HwgA6rLQL9vMJ0ib56sOWjRQ9cmrTiWH/yri6HLHnEovnU+NyAw2o+MjiFWNOotzJMTjLq5Xr
o2Ke5vy/jziElw4VZ+dPwVWh26WV9y3KYEYCBN91tMlFEgwxThG1smZndgNBW9WBCvLJKtT38iJS
1ZrMEs1rR8n3iphIIxYCD21TWGn/Yh5nFeGiuBOBgQU0XrxFwl++p6ZLV98HxblPsx25jOaJF08v
ykQEPdA1SjZyufz5SjVWpq9metLLDFDOmXfb7ZrSbqfibHUbP+p/SNe0wqxe7NrHcv7b20wXxdEZ
jgj3GUhPsbfUAwzIiF+xXyXHb35rXkfxhuWMzRr1VfCv7o7U8EW6VwEGghg8HpFOFfuK3SsTBLlY
41rsK4kbEahZuJZXCPzUKKaMADEEWv9tWCK/EZOS5ZbwHeVcwq7W5Zg92kTiELJNE4vL0uIHIiiU
XIQim8ppUa3Yi1I1t+J6/dirAPQi9OJ6N0JClhtxUmcwRRV+C2WxDD3ZXoRkTB08qCkqJ2GpXHd2
6pQuyDYhKqRSCU9VZ6hUxxTWPtDdvwjyEXj/OkYuSoJFuLZFJCJ+JmYH8oGTfTpyeFieEBQ/sWor
TXtxUGZiFt2Vjq4z0dPGWw5Y53l0a62/u3zYbbU+mQemJTB/pKJMjgHqZjAWtVOBzSObWiYe4AKe
ZqkwunpP8rs3wOWOqyGlzwN5P+CYSHHelwtnNc42iCO5QwaPaZJknwdJPQRKFT2M22TqKk/wO/kC
GUOaO2okh9zUj1u7I2EEQlv+zQklAs7A9KpQWXhnfiOn0NoOeoMUgaF6QftkR24xNBm26Wvete1q
QaQLpF75RC6RdjkkuhOaFTgepe4RlvEcEo14zC3x0SD1HZp6qdS7sjjlTW8i+37ni6avZe4k0nN8
I4jRBe+ybVOTCwGyB4FQATfCWP2cutLIAYMaIgn7RRvvtwFCFY3yLvyHoWx+lJwJ7vkUFR7kX2Vb
Adj92AV1WJQZtof7Aqw+xliYoeFQeiRNAND+FSmDnzVcYMlKF0ZU/YRNgGn6e77QxpkD4DiXtnnr
fB+MObARNiiTxbLlhrsteA6pTONZRSiGZTPla4xSsgax71Q71GVwZi7snATt9I9qCT6XKhe+KNyF
HP5mfhBlvFTFzGApixVocI+W8cgyzSCpJjldWLNkD5Eu8YupIkPqO4oAHG5pA2vy50m/K+mmG1um
ET/3F+CTdtkcLxn5jgfWEve3yoXGp//M4HESqbq0N01m7XrdZdDENlK0UL5dO3X+7Zn61Zes8DN7
PswY9p2nVU/wqGFjRiwaFF0avvy1gGoSUp9l1QlGb0TWVYE/YtbejUgwrrmLJpGnuhufvDeqAU3A
iGsplOH7hMjvx2T6BAbmGW0aRHHjLvg33yWUTv282ePVxrfVWYfZGm2aWCILnbtsRWlrEE8VzzMi
uAx9dL9gVd1OVOVjhusMpa2u77dAcwlNmYvDPNayP628ImFbCfAbM7Q5Io0Kh6yVTL0IUE+v3qWW
iGMPnrRmcCA2ZIrzvXQ4UtKTnGy9s0fWjiHSMGYchVjZA36UzTqUBrsGDMJnxk9I7j8iPTmvDzI0
H6mToQRTexQC1FYe9PZpvefTsSL/Wbt5wZsB369QXvNXFac6MCdkW0wzjXZdwk1y/mLYJbUf4bTj
wZLg1Ys4iJUPgIkt4noddDz2hQqUnnWyx7m6+3/bJL+08YGAVECBaWybGAoK+ci5IcirIxrQI0Id
VuZYuxlEVNM5ZlOC3CGRogghvfItk/ENnQwCy3DYQuUFolmRCJS6d2AfbHWcNErNugVd2M7g+YVW
dtMcyOhwKGf4ovaCqf9MKOdsojmWCNPbMtz5gkePnOfx5H5TsJ3lFo1x7gKLiNYCvcigXB6e6Od4
XmmXKmnYA+wG8Ks+uJPvCTO6xiXNPX19dtM2iSwonrlo36XHZQ8QL6HmXpssiDrv571POlZSdJ2p
UrZdTjPa2F7m5zNfpOhWpzV34aucjdmLp+AqoCGqY99lZ83WSnztju2ThllSdXkAPYnEF6fmPp5Q
dVLHeszYpMqLVVcl9C71FlXYvNhcg1+cTDKl2awMSNX2H3ev2WZsLplhDfuYMLB+0LrIJMcCjsLE
AmRBv4tO3ipuNmGb0uoDoJr1tjjLJfnmzXN5sHrzO4J2t/07p8WN6Eh8ot9hjrjnGTIobwUwVU/k
t2lXAHEZ21dsKwIyMBzju75xkILzie0RA9Gu7A6OcCGBDhBYXhsbF1WnJ0vX2tWT9tG6QC1tBNCC
U4XHDysNepdNNUORESAgmG0rxOXBMVT5DYu8x+gdiev8MENZLgSAjKvs2nUROZu8DBTFun3RoMTk
0ryJ6vl7TQc6U2r9ZUe751A2UNjXCH9A/AA2GBxjE0ZwF+tCON39irCbhZoJQgDopHP+8sq2Ypoe
GMlU3j7fYHu696KINGTHkK2tEWQuzyaQB1nARi64OU45trVPZvovwQZSwW7beFz1JjmzjUqKSVeo
dkz0lK6ItfTBwCCnVp0mRzq4wNCqmbkePTak5AWmfhCUzWD+Z5n2BFDLvObTDccBNTAHJs++cjC3
qv84cfbkZNfrbbxkUGsSBdd6w+/DSkoPc7nVHsD0pi9vj4LpF4NuH7Pfta0HBrIrpZfseqGj+7wz
QeeEVijqxCTjf5zYYx85oNNa08mIYi8hJ9a2u692zZT8ubUrnvtkoe+ZiiQh0MHbLohJWw+B75U9
WwsxohGj15jbUM+jdFlH/+i/na/NOC+Os6aBuRfIkoBbHbv97i3qrqlnql8J2oc2aq98VLRnutC4
82menxKXfDb/hZemEecQ6hzbuD7k9z+l05FIPlaCcj9VAhwRcCAm4Wr4H9iMoh7SLuYtqltnTQVs
5Uf/3S3ihAWU9M8fsbA6U8uAu4sDJrnyZ/GKvKIV9seQM0ZqE8sFV9e/FOh0g5QrlEph1/9/ziDh
kcS0oqXGNq8v1B+CDNTX5XInEsN/aNfkzZoXo1QHYYmdZ3mi1lE/MsWME19Ap3Hk6Q54b9bYIahJ
GHlu9nIT6+B4dSYp5y6SQf0/b1yc7VXMFvL+Vn2dGtkk/OFYSfpqqdTNpJISBS8+peZnf3yWTTsh
ZETxl9VI2Whg5AhrEf+4NwDEboVX0JuEGKVXlKHiWiMp3g8vBkS4dz02YqVEr/C6TNFsQL/D/31R
GXgmsiH/QBpqO3qzXzeyNm1UpNfz2xPtY5fgQKGouZP4W9Ks329s4ax6UKoMijhZYEHlRIbQZcxK
w9mQEPd3w42CgHEwULjhOxKyZLAm/zi1IVXnbijK+qW3NW6hiBoVWfDuoMdIFqA1eo8aqf8PCwBM
F2HQlZjx0vjZ3q3OIKS9BAh9VdRU7gdSoTUgMi0OmZGUk+OeNCCYjJuGxa+ra5BGXalPhbmkgkz7
0W8KCcNFSLxeS9ieHPcFdmvIvUZQSJQK7wzFo3H2mOSYcG3A8t+RiJ65Ymp1o15mAyyyEuuDsoIb
gcwxr7a/E8vVmvU1veourPTcKf+AcXVuY9k3KX9bfrxa1HyRkYzhJjKLTrXoKegmb1WTjyT1NwUS
9O8MA6VwhSmp+kVd5Y/MR6M9tWlL9vCu7tzj8rYqjWHri3bKqZeGuPx2sKcSq5FVprECsXLA98MW
/IOXkEGXlM9Dk2eTcPkY52OqedRvIdmd8g2re+feEYWxwcn1ycxou3rZR55s26kXJkdic6nwrKss
bF0DntnvicVFJuR4os5hYIEwZSVibU559RFP0JG33HeQNCiUPRiE27PP9y0JhX3lBxXAeS+Kpzo/
U+vi8KkQ3L8bn6QjlkWkFE+waWwfaDhVKi4KwITmvOw0NrBHODXbRYZApdyyt7PGGNMHfAaeGkv6
nAK1P+acu3/To21+vQeQ1Foyr+1G1y7t0Fx6jfeHkIWYsRJpvkQpFa/qkiR3vDRawvJk+AMAgyhd
LgQnC2hv4s9BIjI2+pD1+GVQ2/vXKi0AxRo6/plLDi5YoiMe5BZppfoHyLo0dIltUgSdQG1oM9G+
YCoESnx3Bo1Cv8p2pcHLl5BOXEIn4o6s0ZTRuMU2iHe8AThyD9KqWiboiHW5FGZ3TcGpslVlntvX
ZQw/4L36qtPNLSVauDkSSq2WChvUbLGLUTUp5x8IA3iFMLYI6S2bZ7zUOTSur9blZuBsTrmolj7s
rvzz/MitNNeQxfXfGE2OtH4Vye1ECd7U+FmxKO/8sNiDSqoAqERb1ynqMV3fAsCyTWbkg2Woq7ul
+bPU9cIqPYPrq7wGvln2aJ89O12NdHmNpNMCUuyxlDVc6RERnJuRfEqvsHjEzNDRSa1oHkziZLbc
dUpZYTmQNu4r2xpfP5NPzxzWNwkb2bxfISR3iqMbOCmI2QbpMiujf0T5VEHxy/EF982vo9PMmygq
PHHre1RcXf1KgngxlBFvEeSFSLOY6ZzSb2g0LHUgU6OiwBaFHfxTkZ04YxAqEgdj1V/8H8VI4keH
NFPMEF+APlOAkQP8In+0zoYeQkr3ZU87MjXck9VlBfRbNsEi6Vb++VZRlIsZxBGzSc5zNZMakYfK
1fD/XLqQaKjqEj7UOgLzJlZJwTfXg8bigjmmEueIe2hlp635z7dGElFfrvPgPKpw+NwYYkewb/KL
OrrFCnXVeYdlof1vk9hU8v7KEcq5M+bO0f1BAT4gm9+tvto0mWL5xPqIqQzoC9K96whklpmy8eS5
xfn0Er/nZdVg6MC9IA1cE1UStfKDDit5EStQHN82Mc8MpS2tBZTpiyjpm6EfkmXu46IVq2n2r20Q
6GIL01Wr5XYBbcauTVDcZLtjJjjZcYz+Ts6mybuvfuhmnMKMQHqLt03EhDvwNlUMMwZNau92P/IU
Ls1g5T+97hLILtstKbdAf3tlikIhia8uqMTTV7QhMWK37MSretLiFpC3B2zqK4PC4CGCTLkGR4C9
wzYgAw1+I8ipDHzAAje3m+2Mh+IPtxaypEMl+eIFnzGf6wEmhTp2qLKWgCMkaP/OHrHCDyCJ16WR
CRHJm55LiZ1TM13Zw+373Y5RreQqKYyYbgmM/+xCC6sfmG4QxJgmASTdCvaD59eWBt3LfnqLOKfD
RUedONegWC9L3UaD7W8I/mKambiDhMKpB/yuTcxJcCMSuM4Lvyfj2v5EsYZn1XbJq0JT7G0fuqYx
Tpxi6rgrGeAn+CsaChsMZwIgrK8BTOYZxhyfHzyjQSoaG6O6h4sKbTOe9LSr7t3RK5DPKUlzrKtJ
UqmUoK6DKeC8iBoIc0ymsrNdVRzRGlfdr5lXI1Gb+C9+6FFytSsZAuvNybME9jRaLHoFqeK9xGbC
kjZnXoPKWneZp/1FG3df90OZOcKrYUFv3I2rMBJgpur3Qg4vmG5nVLOcJtdhvMj1EkRLD0dEFlQ7
63Ltpifb6lZf6whsAbiSgDqnNOurbssnyn241X9gzFTGj+RxuzLBRIVw8Tfn1etu2nVeU0UHV1r5
K9vfE2fcsV5DIhCNkxaM9WQGP8hjky0ev6C+bm8zM+Qjdut1W/g4jrd3EwJlqPqqLjxqqgJu1BfI
1ztLfJdxyRhFIvn63lzyWtEVgqrpThYmugO4rePBO9EEqrRaWD5OLqyHSrxy84Mz00ZkRQl4s9Ts
CX5bGkPRDG5qHqOUFZdMeLcDVuOq06Otb6uxbiFG8bwc0g+ELcS2+wPpQPMSzpkDuLomQz85NxHJ
xav4k5OjCkRRksbDwNVz11MzVE5caWecfasAqtGTfEdK23qzlRv7J1AF2RyNkgI3x9XUgzn8KH9m
Uzlu/8dklR75b17GVsMn8FR+R4gkFLiF0YGkdDdZjtqko8iQ7TYVG0WD1zbjRHi1Y+b26F+DzOCZ
TywZS1Crs1v+ZiWKnzMEk8d9ZuiqkzGThmcE6BWMItQLtsk2tsrpvlcN/DDAI1Ls375HEsrEHmsn
ChUKjooTV2s7qB5jgFi09G0gg3JubBS0clGIJ2hU1Xunh33Oond5Xex4+PzSrlo3JIgC9+SPST+I
hVcfPWG59YOSnoJvpWFpDYN3SvFOdboEVZKXNtWPj/47B+nfg02b4XQs9m0539Hcb2Jz2MMFUveo
7FsbBaq91K2W/n1msQL28xDdmTsGyFZXB3hJ/wBRWLH/pWnfk2yg0WBgEn+UA3UR0vtBY3Q/VsKj
G6Et8xSkhqrIzypfJDQ415RiEAgu+4itsSaLLvgorPt1RrUVqitqkCZPI6ElRgElvRbBWWUnyiGK
pH4ominDziws9RynDhPTxafU1Ed+dT19tNj2Hjni9Ty68qqvpG1J4yaURFO18EfnOMlprdyOlYed
ReZLaSFIk7BvcLsZ2HDCgBCh8DzK/EURfp/nIA5HVWD1zBc4H1M3eT+RF7APCVhNKqeySgLPU3Ge
z04skQuEhEnSvoZ7se/eIiAdLjTmZL8JTE+KjXCz91gUL8kAjuvLpFPUpqy2+wTJA1E4PpsCJEOY
pPlMNFTGaGkwNqTDe3ayO3eBWpyF8F5jR4KcfYs93YyrjW8rz/m52wb7i1WarN6GWSIPGhkoQdQ7
QnSrLjs7pBQIdQZewRNreZ8YFD1RIJzyNC8bgBAyW9lGaILMf3tJV5EU1DzRdxyePnQB23DJ0Uex
H7qdmBvw75nf/IeZBx9BUOYyaGg8PWlEj6LmgTTKbXiCVsCYpWtpvzDEQshm1tYc0VNdjb/I8Icq
mzBWzp7qSaxTV+EgZbOP4UpaVRyMfGv1g1wFS4dPeTSp7HYMgaRXdQuafKRywU1BrRKyTw+7gQzU
siqV5KdaFLMekHTz/P9nZW64xh3oUSl96u/185bMc6wo74BgAZ4eEmqMbD0QSPxBEbmO/9mxx8r2
vDRdrPyT9YSR1/JSdbqVC9yO4BhB88OtYx0qorqc4S1ZpQO7e7rFJiYz7/PtLFzBmfNk2MoSnghy
6A==
`protect end_protected
