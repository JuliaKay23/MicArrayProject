// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
A40hYsHvrgyWaZFWC4Gzfw3UL494bKJyBgKPuJNE1+9+9FQ8olbU0VwGW39CTgQbR6kiiKLfOugm
PdlAddC1HUyemVOetAj8Ecm5dyegxSSskooD0X7mynTf4KQQFpF5xPeEcpxzIJbib9G5a5ogRuZw
TY2zluh25wF9fEpccS1stJ77DTJTcMUnYECPje8AuYe0SbD5iczz2BQizq7l0ItUV7HIqgjRYXTV
i7JpMRwYp3tPvKikLtvHqolGNYwIFBOkG216oIdTqW3zc7ZMusPEMRkpIa4hsdzU7V2tkLGZ2SD1
MjWYny35MVRUTtVBGBGR3Z1Iisj0h7SqLUuVbA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9008)
mTy8vanGWesCnL29QCre1FfJR2e5iGmFubrBvc23u2+YSkBrf31hEsDRyBMs/ocRIQndf1sr+CrV
Mi1Mjm7gc++uSn5q2DAkUugyZ8LE7MNv1YOoajl07SK1AcgLO2JimASGj489qVfJq9rJ+AyFcqYx
9eG9THb62fUy12aKon5MosKQrl/tqj2t0qfBWgmIOwrqopEUdEZO7GPHV8dNC8CLFphD0/lGqZkc
B11foltL9ogL50NDS4a2LYYuSHcnTfCvpBdGjuY733t96UrNp2/eMwrPDSu4w9eN/BFt15VZOtOu
WkN0TlDPmQDKGBQ66GSGH4YxMFrqLXHhrvu8Kh9onYyazIJCv0t9dTrPneSeYxx54vHTbQIHlluF
qctnviA22v69dLputvtFfpJSu9kxdL46pjWtuuDH8JHSTGwwVcyN9gB0l72Il6pJO3jHxY85eclK
/iYYgMuZM5MEb+s61c69IAWK7/AyyILYwbDTtq1PfuECbbhQJ/MgDP5FBl5U1fZ4EUEg1ZPMPmsh
C19Q0+7Xi9ocSpF55L+NQw5Wk0LsWkJfjj011z/BKJWaW0HG4R1GOmBNwCOKnP2cw93XBHYwt4qJ
69jbTGyV1i/ACoGfMR6vx6bGiTlwqkwQkcoGL7lCW99nFKNVLxXPHri2muUE0mKjB59W2FsNCbKc
R3u8yt87B1+bhtVMpnUCXxzkGcU936d26RVwjiREismdf3nt65oHJKMj9o6jQSpeyZIRm2uicuuB
Hws8ElnPRyrKXoyEH1vCuVgF2O/GmpuJirpp0aPdwr/1Qhwqvz8hErwbUd/0+F8BnckXcqQ/6+LI
PEsGAJnypBpp+y8rHPDLp/XXMqsjV6dWZMlsXu0kAV4yJutSGhu1KNcDm3Pf5zq4bMEBqRZcDqVO
eplOyLcruGOjcU/tuuoZZRrHAuq3gWe2mrbqz27TSJIPKpSgHcUP5wqXFAAqMmuLZ++bPUcdwVAx
uzC7xOcfwWMaYUHcGgyvphU/IJl6dfYaE+PPh+LrPntvjHlndsa9L846TOrjw5ri8JxQYHrHu3wc
tUaqGau+vOIVs8gNJHYTZGduxVg5KrVqZR3qfip3WlQwkY58DamwPvRbEYITqG61eAH/aARRQLMx
10ix2ui7saS/viw19RUerc1PUMKAKzE2Cf6xfly5Co/gxSxq8LLSOPu5uhZj4BiXBwklBUOszFb8
i5AtQnv3vIk34TAFUX936jvDfPH+VahdVBOuqGqHtxfB68H0sV1/P6S66rwUa9eWYAQCPZXlMQcY
rasNuV+/2eEdExaDMCZDHLE6SrqYzu5vhYdI+wYG6sRW7F5LFCNNCoweOtElk8KXCkNGBss5LjoR
7y8AxhL2Lqm2B1AQtPI2aYmBq9L+JcPfMogN6Bva4CHee70MJDTxex/RlyEOKZ0/KWz9+Wy07BqV
tL7bYd/ymQg2H39qV+I4/Jeopyw//Y8Sc6CDr2xViElHCkHr1GBVrsG94YSmbSBsTBeUsTXVKX46
iSNSDMBg35S02MAza83XXRVpHcXoWZtJAJAjcaz2cgDcz7HBTqgF6DVEuBCa+jqPE+QWEHE00h57
vn6sjfeX4TQUSIwPWT+fxeAlloGy7hNEUYTaNAFDiTIC1+eitfMfd9MAvoKORvI9F0mYD3rIbEzQ
dpBkvh97zdloA1xfFKIbnpVGgBW6oapLiChQFChC8KIon3UpDUfEFki/dtSU5MTK0bwizl4lFbDu
t5WpmckP+g+4XzHSlAPSJ40QDWmRO4MeC/WxUGQvW1nLDcTIheckQ6I/CLyuOQ6BLBaVs2sU/eKl
ar3FTOSbWl8kwnkb3CPtNZVtjijhKWQSMEzwDRxhmd99mA9iP+k6L5Y23Ak6oUHuWEqzARHcjnbY
on7LDW1IPiH+AzuR8zB77EzDhc2i1Hrmd4cJ04af2o0XF9dtxtYS1C/T713sCOgEafR70zmrLBdy
JLlVkVphgs9GSIVOQZ8UBs419XrlcD9t+PgzMiTEDqsIU4vw3wrc5f3FXW68bfCkIVL0MNM47Heo
PxhnndPbGLQmWQhwFzkK8q/8DaN5akBF9Hmi1hyoaIUDeVZT9DgBcWvQdZDkc4jL6lD4GbaPL0B/
As/TTxE1t9Vs/W620rfOekkNh9FPTghzcZcSeTZtmgGJFaosO5b83RITtRxQqEUotaEngvPKor+d
ZN9fDbZFrTrUpsb0YkutP/8LpR+Eogtgm+xpVLwb99L+MS0aN5IviaxsvRoRufbi7jyCf1uCKjIT
hmCFF0HTxkbM2hkYwWADo2uZTnwpUS4/XpM5lc9qCOVKtZ7KPJeR8IXqAngz+YXRiseotwepRnhW
gbPxOOEtSKl0IKGj5KldaPVEsR77o31ePVPuPeehZQBW9QUHYpmU7avGZ3wkpd+1c4IfRHlvlEl5
IyCFWUV7DnbC+VRG73Tay+9dJUo0OzdyRNGg0mNW1wulqAJE3PiyhCfsH3yHIhKpxJreJ3rhVZQe
fV8HxK1YtXa4zf5u3ECELRotjMuCEfOAOJokNADtosSQ/N6WEMAwbhVx4UxKn5DuOHgXmk820Vkr
1Mr9P7jh7xAYKeusB4/N66IU3rYTfRgKwSEPPomNBbMBTUS/GDqacbdeB79WfJVDpNR177FJ1olE
kw2O7ChQ/baqc/mOsgm4dRmxUN5CZUAWFzWYo18zY9yCORk+iToNgRSUFOXIPbT0Zxs42XXT8Vy6
h3R6ECsSNOJ7h921CUC6Vj7kiP7mActzAJ2kw0cbYeIgv21PhX0p5z7ETz1L8ZOjnj5YNrxUzzup
sj4PJqL8MJuaGzKeww8Q5Ym6VDRI1nHkOPbC1CtiQYFpy4lkexiJL10kkXAj5xSuGyI2VsThLxNS
6G9Sakpb5cdJLiP6lcEhyF4jOhEu6/pMiy+AIT6mJk9/mT2UtAR33wEJOLxezxAXYjfb0lVYWzUe
3zGli78H+gg5jt1Rysb7vU++J9dcA6RTil3w6jyZJnGMFaeavjywqsyOOaQNg/1OJOOepUJ+F9ud
s3cqjhirir6RE7xLA+bzJAG5F1ns4Fr+S38jOmktWkZrfhnbYbSq4/Fcqnd2f/21moLAy+aqwkSI
YS0trXnUIfI04tzsphMzS5DBNsp8LuBE+pBF376MTpbhlSDK534maPE01LCTu/C5anW3QZYuZ22e
LmnxP/7vkc3JC3/ImUo9iuRnOy0tDe87+lxl53dc0q1do1UrbNo/jPLjWy92BG6rT6Brc9htOA7o
/uxXI2pb8Vo6wneXjtbPCCQW+3u+ly3T//7AoJq5RmtENhK/z81E1UOEOw7qvIkOpc4qyT0DMC1R
uzpa2kyxPz6cej/UZ19DqASynLq+0QXyrulc9/0yrX9SiwO1A1DgQUDnedrhpZ7+5n0kQcm74FIu
PqhzNUEpu8xNeiqJMNXPJzaxPF9vixQNCI/eDtzA12pWZ21nG8ccXk1wFLNBazjg7lv3ewWjtNE9
BfA1Xzz0YbZJsz1ykLkvMISzDQrv/8ythEWCx/g4pNRYoPCtm83UzLmJPmBAqm9ceArnYOTj6hm+
WdSZhpnvjkftu358XCMrT8JoeTfKXV2XbS31kaZpfAQ+82R8sdhPjlhuVQj4YcYd+mC9RsbinDjo
AjA44fGlgqdfeliCYEyuBvoB8EXDUv95tlvWoD3z2cIkakXnvlJpP0h0OdRsBoO23ttMzPBjM3Vj
GqIdMZHbhBYOj25BHBoLXv8cmTUW/VkzXN7VTVUkbM1uMGTJDNDPX7wldCbsh6BEqIB84opzsHW5
MkRzUdpAci3PsZ9MowBkGkNt4y8OF4r/3vHVwbr0wEmOWWMYYY0YY2T3qCKbpHWYqS6RuB5NbqrE
9TGEcgE+r4Soe+bJH8dEf43dZampPs7sX2eR2p31mvkYpouOBJA+Y626tWxnIFlhoXcd7RPwjT2U
AOXgtEUHnmopTQVkZqn4TP13Y1XBKmPXfzP7QS7A+Yx3JXIOGKLhPRAoIz3KWnoUFjO67WNkLmm3
Kpa4fRip2k6tmUaUpIeKUjWwmYJelG9hPKEspQT7nMYXaR3R++ow29kTq2aJMvVBmSjVQ4LQYghe
fF/FKKyc7C8duWFEQBgvUyFSQFuLYyxmnHvV/Ec0+TU7tuoowfLdvCr8yW3rWpL1oX+lTaLSrIHm
l5AVTqDwXDqeXzi0rZEV9dzCDVCJf4l5tb4aT+9u+IxFl6hHdWcq0F9kUYh146nHdYtve+TGF+Ep
J4vXTzf4fovf7i4IHuY57FKlmBPQjHiM+hiZcHCjbPdd5eicp9h7UkXF/zGfqH9zl+D87PDRn2V6
Ia4FjISnEo35ZPSX3uT+kQNJCDJQ9sSctujwER9kiZ7eQo2mWScjvMQhzyMdTqUe+mxKcbBL1DVh
QwWzeRmXwdP7Y45yB1EukkqTyTlPH6JkaUqM9fKoAvQ2I4EZQxVhunWpKgvCXoJMc2/l/PXQQIU5
UVkeic4SyG3L8HB6zMr3BHA/AhA0l3HP7XZDixDIaHZQvlVrDLFA31hk++seVuFZxVVqmaAZ4+lL
FZX19zdeELxLpNkCrVxcdtahJV50DTsH4FoinukcVk35uGR9BYzWCHapkYIPbYtVLCLVT2Muj0Op
RkUhGavjaRnRanhdTG5UKMmS0GtnUIKY1BHTPuhIQaioD11ezarco4o+pNGu0d2g/TmkIOAe/Zup
TANC/Kk/ny/KglJ65lLn00ManSyFP4S2dNyI4/4cyaE50Kcjgcjpmb2iOR5pRfsrCiX534JaBGjx
DbNdql6hOgG2H77QopS0tItlDtQBj4S1WCOFmn09KvEKzgRDGi1A84VXX6DqBZmCqP4Ovo+YZEkn
RIDbYpvZMAAxMP9FXmgQ7R+beaZF+YT3RQG7BTHY1sZXeTaxpSbKVv/kHPCSmnsVfTabboIJG4Ry
4atZGtg2/1phwUvUogyaK117aPSWuQVo6JpGEKju3eubX+PuJCatHdy6/u5qwaizPmCPsLLw1HkP
xP2EccD8j0Y/wSPC2wvfjub5P2SrytFb2rdE9BfsXmG6+OY4wmUf51BR6MpLVWQWGLTtU7CBAtNF
VNgVCDxMWgylKEd862ut/4qlkouusU7jgMZFFqJrIUMsYFKLWvKpboaFPHezS6oxjulNperpEW2p
1/F4wu0TdymeSORbHScX1B3Dq9RXIhacHkpBqPuCtpWY4HjOjjFYZEn2sDQn2nm74PdOl1Laeovy
uAGbaSL2ijw4U20EKflvpFWR1kUzSA/++9isUF0pVtrHLRKmmQBH2HNvIQ+e7y3zPSDTipRK76a8
Rw1dsn6QKPEO4BtrmQ7NgcUSOHh3SfiktjT6jHRys4YKOgBKol8/YZfKdGMuGfnuS2oLKhiThWKP
4BNgaHB4NXDaNDTrezdaX2ZEhYyr9fX5fS0fNDNLM9IeVKVwqcgM25u22b2LR2p3ZXHZ8/UclCxg
7S56nnfwLJI0ZptTxwLcL4tRAXfZBPv+wAzNVHq/x1WaJSizPELN8LBk0ceL+wdm2F9vY6f49gEo
hnc7gPg5YmUL/BIIMwV0TyHUhH55/0TtvbG3ZHXEbAJxJEkj2q6MmZ3yPmvGkHmxdMGxRy1KSJ2y
6g0X+Ls0z1yjTankeFjo8sKMkamWKX9c35ZKsuY9T6NRNs/8Kzw8r9Gt+MELw4B7PX2urlXIC0Jp
BdcKs+Y/A8vL6WI1NwSzFGYpthzPXdl9pR0jxwpg0v1S/QuoFeQVT8TMXJYRyaSrdHLdqyEhvyDX
x2Q8UHeWd2UA5anDOnnLs7OLlkowud+ByckqgJosAbQG6A+rR+ZQJMoP2XHpQOgbD8a5YSS44Uei
cpB/WrNgL09c8Sxe1oWGw9TkCIhfitgLKFQ5hqOIIi+XIZu3UK3UOD47wzjMQyL8Uar55v+GBRuZ
wl0cpLU5kdGiUe1iW/JSMkq8deAzFr+zLRt/iFRrYkaiqmJ43PpsAaASdsgfbDQJeYicnYGUBvLC
6UcXUdqb6vGbvT3vBZc6hk9yNU6yfJ/I799fDL4pHPvOnVgQiyuCjzKQiBwLqJY+nV3ue0WZUBs7
G0vEjupnLK8JOvC0FttZV2vM/XQZXSv/UgSBstC+yPhdng9FtVxKjZcl9fHu5guPkdYQsFqBwaeS
wW1bb3ukUTR22GWK7Zks2JGt3C4TMBOaqFTU1QvOkl1/xjlhnMGE4sfLwHtgSYubtOVP8rxAIjnN
iFsJWuUbZxc46QXg8CO74Pif+4CXIWmGPiFVJENd9gKk+rEDYBeRHomns02Q2zQ+AyW0l+pNYa6P
AjuxG2nuLoJEd+GnGpXM5JbQA55EoRoRrpHVYNZNGXfsPHFNF2jm4L0sCMt4P83uSUSH2lr2BfB8
1tXfbcDMrZAioXML+QifmzyQxo8dBr8Ek9/SEGO1pBDiRyLyyXI9Q+vzuaIpCnf7FRbG3r3o4n/U
CzCV+Rc1hlEcsOwpfzh81MRWUmt2KGlsbPHWlNY+0j5KQgb0FaotVsQDWlPZOiklaSd0FmMY+55w
GePbV1LowsbRV9OwLNTn4NjuK618Tvgq7d+BTv9+H/xDbG0yBTwnpBaUD4Tn5DYjD0HIlUm6X828
XORkRXfk6ldEUgGi8z1ZW1IwZx638RbNBYYlEYwK+r110Nvbj3fs8i0Uth2cCqFXLbkIKPg57NwV
3oXCJxLej5+3EHeHCYifcO32TZWMLHsOaoOCigGTrtMJ0Op5oZYIJI6H1EYZkq2aHMPKyLI0480Q
3ZYR1bv1ouS0hINEiA52k4rS86BgV4ahd5Q4d19xhFSRzj9eAmy0EDQYGBrSo1K4Sy3flRZ1Pu8F
imocwYda4MqeCkF7keRVbxLqREn6NNTfUlwJNIRS8CghBX0kDcxAQ/FRE+BiYqYam/ajfXq3WYo4
f9kF4BkdXSMxn2VhlRJguBqLUNb/EJEE6gFhUgbdI8MYHGs8SbknaMiG1Xz7OZR4680qOMSGuhka
nNZg5i9tRl9w1LoM2EL4m+CcApfZQW3tU8rcKfkshDcnCA2oES1yzeDywiMBae/3mfyziTm+g4M8
QJItz14Gxy93e14D3gKUyw5IV2KvLfoTdnchRUuHxfaywOl0GQljScGNRYY92Y9wpgUkxlwKjyxg
IxSaQfoj6ojoWcii5XQRgnDsIqpsTWeP5XlVzRJGAKPqqDItSbKgtNn65wmcZerYnCf6O7xSAung
eKABjk8AtVw+CvnHd1JhSXXVNjSdf+mjzomLFFK4pt3YHsuKHSfYCrZRVIbtWD5wMyaVvBJ12YNL
/zCP3GJFdLnsZMQIr/aVd9ffR87qPV0X7CJYp2xX98Hc5lk3W3DyGLIlwvBImHelAZjwy3T2TNZ2
BYtiu9I32e3sijaUcDFZkmbH3kn6biLgJVfYxIWjrLr8YoFJG4n5Xx9xShYiS01iR5/dVkr49b/Q
iJfR3S5fQWqBP1yM7UJG3nsWnUN3yZHKRJUyY9Im8ohQNiSxKwK0lEN2v4Lu9hgqvDsbTm4P09+G
ew92W3k4jeS1lHGQBUFGphzH6wS7AhuSCKRglzsXhPdpvSrhH8W3ocWI7TX2QXfZ9Fqe5CF2/r/J
YWyiZCAYbwf5XQdGHsZpnQFfvZ1oobCg/fipQ5I0HhToCwmY1Mgj2HTM0ahHUfAHZtEUv8MEpPvG
mik8AclRNv+KXWS/QjghMuPkOHvstF0SelYDtDnYodaNgrM8Zt7FvtTj2ko4OWM4+rG8OMgibGc5
WW4rUMehcFSjkEQrUZmRRCN10sG2R9Yf65e/FFYM/UK6DhLWrSRHecOk6brUt+QsxAmrTFBULWW0
W8r6qJDJTPX9Cnhw0lnzQG4NvYNl8UUgMl+w+kR+6jpA9LSd6DGjjHMs3NDEn2Tqn3SN5YJb6LRN
EcqRzZjxJX/6x8HaOVbeTA5vV7009PuqINmd0lHWDCZYQ/b6bkq0glDo8QrRKxQYyxKfR8TWlfyX
sCIarIYZn/gFqOH44oEOqfr//VUnQmiJQgPkI3rlOueCJ7143EG/m3JKi7h93AUZYEySi7GD2hzm
A5Hjs52mS6O7V9faEQ54HawRB6/pqgipQUzXfi7T3lLnGeFEJPoR/ZvE8LtNppLqBt5lxw7SX+XR
i9YMrS50qj3YPTIf1N6iUsCcesIAwNNeil++hwmG3dckprMhXlFx3nDYqODtogUNxcSmkLMQGhHn
QKo6z6qcSiU3nG3V0SzV1aHYucHVs54phjLdMXdDjszWffFe3FwRHA5dWqqCC+J3+BQv2UPKgt3/
tvQyh8SjqySh150xLJaliLEODbN5ArroPW0eE+N6nZQKy2Vj8PbQUSAeT4+yCBgsULNF/12F7jgf
Y8PlnD/PdJufR17D7zOfFi5fWJ6jtOuiUGsdEEFC7aeiOCOIiL0B4/5M8vjGeT1aynelGY6ZNxkw
Vbk3eNE4u6eK5aCOAJGlnesfwBrRm0QhdIX46wShp25zZv04PJQEV2JjDpog869HhHd78UsYLvxw
fyTqj6c5kGCGWrR1odUnhOc/nlYjxwwVaCP7/ERzdPCn5aB4T+kOiq7WOpMEpCTfTH6LY497HG7B
FseSOFloX7OwRBM+rXfEqU1gpOeZenlaZnggieYykHjjsZAypORBCEGG38FTr/7QWdOj0p0MJVKO
QwKBCKASUW3DL/zqjlu7VRVVFfhvZCwsDmrNDyTUkVQrR1TdIeFJzypTozONFOD0HsbstX1BGt/z
8UzFNUhsmjvj2ZMD/q66D5Bienw8DNzBwEnHaASUcilu2Jv0GS+Ax0NZ9IAdLNiJ+tTUiiebGfWm
MplHlILheuyTAMLxf+EKemooROsLps+hUUJCLNnsl6qSUkPpK+cw7RcH4TQ59NvtWwVI9caGPG/a
SlagmB0QV1iANP1+9XOqR9RIHp8pWp5Gi112k4Mt7dD/eyNAjL3zgGQC18R9Nq2wRGnQG+Ngh20H
qePsNCbRlR+Fmc0zMIuYMutJKUnRHDj969KXSBv+/8Oo7YAmcWFBXdalCqa9p50TYrEWeK3Pficm
Uhb8fKKMgjnJQ66R2c5LHGqgqm8Nn9uKIYXn7xm4vAWh4drkjcRJcWNaOjoLWxuot/FXZEzxa+iQ
z1gdXgJUg2HBGNCGVBlrZcdTshLaIMa/EyJdjtwpc0v1GL0ZGReG0c95/txX7GZhowQcqQYB8R1y
IAg0XgJkl6jAm8T3DmMv4ypa6R89A2qo8o7MMh3xxE13Nznw3c+L3Qk+obZK+eIsv4iD94/EFZxY
/1YK6O3ZmYNZ2Z/hjcIvQLBK4Pq9GdlNWuLtB0y6PuJf0hrni/zcrAN8gPepwOivAsZii2OKTCOF
nOJ4yslm5wJFCRQwo0lQJSOEjNHNpn5bfIVa4cPEh/8dVD73MDutPTN4st+VF9zjbSI/V0+l2n8C
q6vDCrvhrAlEqoOgtl7Mir1WI6od2s56v0BVB582JeioVi4gR3wyavSb7K5ZuC9M0bw++pI9P02v
tfk/rVWaGKszND1R/Qk9pl6w+6esluQX6oNMvyJ1EPSxa9tLgY112rkhIPzclZ6Pg9UMPmxZg27b
UCaJorHKE3tG9r9YWEtVISxrUl1C7lkyM8EefmZZUN0LVkbL7AJClgomSm+HZvCGGNXvOPnKom+w
T+hZqDF7QiRXmZaU0OiJcXIgkz4bEinvxOqJZVmLNJ9cYAp+iFndZYyBdfY5uCFVOZguYN/VrcQl
tKAtm2YvQfzu10Ar4yirAoJ1Ij7KgGjQa7TjfLGgG2vrIS5uhHkhhbII7Msj3fcJWbmO6WfeezGr
TdhCbTTGM+PV3ZDO7BFh1JTlTXb/te1n3W6HAkwsmOBgq9YagE72AmzSvWtUE2J3fEqOBV6xSmne
RLJxSJkGTTbSjs7Ot/nvU163Z9XAv1CZogGTkEG+2PW3mJoOx8bV07CWjqnRV3+A7s9qXMLYoB7B
dfXkX9IoYwKunCY2Mq+KgyIXukXrOz9SMWmjYGm6zBciOJsWkj+dHkpObwH8wCTvJD/rYVikS0eJ
laQc1N8N6Gb4cpejdgr/4NRGHrHzkQOpGtArCPV5GXUkwEEhmV5fXfBJt2HV0OU5rHVSDtN5L0i3
DHIqfRK0bvIeeH7q4oSrLRmj6oYSZpClTwMIdB6+akZwP1h7XGziXM2a6qRZx3j45eQzmmVnziDK
vNgVhBBH9XUgjWQGDZKxhu0y61ymeipGxR+Aa2SWfbsLaNAyXDYt8BERcfXWBHdyu1Ml8gAxHqnZ
o04RQ2kC6BFbO3gOiQveG83gNI7SYbPaJSfNtQgjsjlcZaFu+npsCccjOKAfFJ+3lVCjEyk6w//j
1Cp6zt6vEFD1xOb/yg0ZNe2prRAxSleqrGDOB4dUM4U8aiBYnDQ3BABcZCZxNVBA/STB4K9Z5xIS
XQ+f0oDeRb1nc5lhHHtrNKMiHgz2pDZZ9/h7eEIpNfcy1Wp7Lnhc00MYgZMat2N4hFJYuIqZMd6A
JN/m3rXkxrcJTZ9H2StpkDEdv8AytIwMijb5pUbuMqt2sl75UGRCD9uEXSc38wrTty7Yz8cdhM4a
/bI51mLOKsKdHnbqHBTn/P7ieHQ1Ta0GT1lMfvEgmrs31dTJMLh0PJXDQNFogTzVCQpNCHN4B/8W
VTwGk83Bz+3AAm5q/fEHH1iYE3hlRLCgTiQo3wJU06pXTmnsKwV6Q/6Vyd8u2BW2PTO2aGebik4c
GMHjVlkqIrxxFT4J868Jwo5fa8yeUswQwii6I/gpSCXFu97Bo+BVWv8XrZNnkC4dadfgIiaf1piR
Y4Ia4O0MR1CE0+W1qT9MHBcl97Hn4yfYNQGL1hNAEXaGHQMv8riyqF85k053M3VcyzapRxvHJjgt
rNa6cFkKKl6NhnlQx6CJkIl8/I2x0P+X/JBuYfEjICfZ0ngaD/4/OPrQCq9XRdWT1SRQ+W8nXqo0
eCLF/9ddcTdaFqyQIDobUyYI0n4N/Te/hekvZcBHR61vOr7fqpRHx2m2mmH7nHRSb0agogAYPpQ9
/cTpUuPYQXoZMaAoTK+tQ0ge/RoPxwLTf8FyHzM+2CpfU+Qud0dJY9S2yW8ELTgjQ9T5+nF3oViO
uZflgezJmnpN66t690glO6Y54WVTcsYwdt4bscPHqdO5Qe28KseKOCpfXkoyIMn+IFCJ3/ZO3Wj5
VN/FFBcBG1qhVj+ODC8U83FpJNEpI9bgreMdCX4gRoVCGDVxYSmF5QB7zL2XqYNi57MBtdg2BwG3
zld0wQBRIWVAM9xF5y0p4l0040CQDbHKuwlfUVskDptGND6F24eUMpoZ81+U/qLFqoxKzsupZFgw
wcLzH9x3LXSQn3OYv2DFtn5FJ3kkOyQD6/Cxa5bb6To/TTdTRO+pBzDOv8EXhoGEC9oxU91YaTvS
bMQdyuVpa202yJ7yL+W7W49SAspsSow2kBzMqKEViTYG91VPi9ZzC90vAVf22xFXoMECin64ei2G
FanUUMKpMuEqqheTuY7howQjYi2uN9nKHAc3AkKVBc6rzVZ8TUG43+GUQyKQeO2iN3dRs00iRaRh
yozcETeQR4NEh7/7Ra7poL7Q1y0vwKd5BHXEMDwffQPgFkrjeFyqcPQ/0r6QYSfjv1+0l4azIotJ
oDfWEke2an5fxzttjtoZhAquJzdxzYuOjkQlPSBGzuiAuzxTCKhkLrntynBmGXmtT5zf4L1cNSQK
hCmhilB8GBWj/3KIncLRuOFB0fDZrEAomISaNbjJIVTYu65F9TBJ/ooEcher36JtLMq0a34UCDIM
ZZ7JqjnjRw/h5c2VyyfV8+nUNArw8/TMZhMM9/BO/I7c0Dx8FvZ2lF/MPRN1tTA4R5jQ4cqOPQWf
pxFGee4mm4CPPvzX0HZA/6FVyTZgRlJWi/8kc+/aGrBQmazl6Drqxj3+cAyszdPaYoN1KqI7dXd4
k0BarvK+yoYs5/MtwooQoTXuUI+s+puoS8d29CvrIeLDp7KH9lhkcIaQx+OT42/JAJgBIzjcJsL8
ScQ=
`pragma protect end_protected
