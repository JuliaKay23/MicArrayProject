��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V{a�p��H����.T}��/���{2WA��b�h�ű ǾPQ#���� G��Y؟� d8�Z��Ut�[��0��yg������70���yF,|Ɂ�/KB�D��)`J���8\��cq̺���������G�sf�_�n�mm­8r�\�&ś�#Oj�n���J�iI�l�#�j�j�����)x��Ju� AϨY1uw���Ϗ;N4��/�E��_O4ʚ�fD����g�lH8q{~�glKi$�A���<��E��O��<
Bl)4��)xe�Ηz���R{�p��N0,�*8��G��Y��[����?"EڙE�G�㐩.W� ~��W�"�`��&���z�O9u�P�d����Wu��st��8��ʪr����G8?t7F�
���!E6�Z��H�2���x�.�r@�c���ݿMt���~ZZ�)�D��j:��&|��g�τ�d��<P�T���G�����7��-��{��8+���L�]�/�|L���Gk�S1�-�1V��;j�4tSxѽg�i 7Ǳ�/�����ɣ�-���wH+s��{>��"z�cd�hڵ/����`�1���.S����'Z�l� X5�Qd�wX�K�ߪm��6
�\�}�е-���s`Wh�����FkCBb����Z;�G�U>�x3lU�d�tg�͹o[�̴FlvL��N�� ��m%�~���,�x��"n��em<k20sFQW�U����Br]�@Ԏ��f{ӳ<d����R�`��?5%׺�����Y������ Oʇ�gp�6�2�|��&z�֎B��]�gb�d4��OZ-��H+��G��$"��"��Ny|������c��=�'!���➢m�cgmD����7$2��we4�4�U£�!����WD���|1�7��|�X�0[$%�����-��cZz?�Hg �=LW<��l��f_Y��3M��ര;[]C4��m�&�����6�����G�I�IQ��tE���d�� ��-�P�8s�}��kq˧̠�j�DS��`]Io4��3�gfu[+���S��.�I���Zʛ.={�Xia���Ok~��	�K��8ڕh��*���:�M��7YܤKT��b-N�-�=�w��������!Cc������s����,�o/RD>�����o�'���������#�����sɃ<����E��O��n6��� ��b�Ε�S���w�����O��ػ����Lm�C#2b��N�;�g2��t;Y״tQ�*���	DkG�j����m��\�9ȫzr�A���I��<�U�����l^0�/.�ݭ�i��SemP��TSd^��z��H���K%���2,H�P�c\Ğԡ�H��t|I�=H���jk��E����*WO�s"�a�'�x�)��'����đ���*����e���@�}�]�V�l�@�>A�c�NgwL�q-��Deъ�I�e�{=e�(�VM�Ks�&�X ���Δ�4�UQ��g�5W�K`f��Ɨ���&�	�����YǏ���V�#�{��]؇�8�;>&��`��%��=A;�r�K.O��yJ�V?�?Y9%i�N���Y�И&�I�f'�Q2С���I�s���ډ�;�+6����|ԋ�J��|�m<�Y�"bϿ���8�o���@��?O�u�o縠 �p��I�Z$f��FI���Z�BR�t
�c�/�"I$ (�1��YԸNt�{y|�j|���H<�@�Q�"d ����7��"�:F��P,�D�C�ƹ{�֋��ˬgĲ�+T��t����,+�s���#E�C�^8��]�����w_!�Q�ӻk�/H$�t	�z���'i^�C��2w���Oi�QV^�8uZ�؉l��gά�o�~�8��R�5)��@�y�S�f��o���#�>�|�soyb���ɧ�Kk,�!Y@%��bo%*����\��2H�:��pD��4�N�(G,)ݘ���Rbr ��0����i��<���Vs0ӑ�)pa�l��0^�c_�p\���w��4o:�l�gt����L��<�p�F�G�