// combined_filter.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module combined_filter (
		input  wire [1:0]  av_st_in_error,  //  av_st_in.error
		input  wire        av_st_in_valid,  //          .valid
		output wire        av_st_in_ready,  //          .ready
		input  wire [1:0]  av_st_in_data,   //          .data
		output wire [15:0] av_st_out_data,  // av_st_out.data
		output wire        av_st_out_valid, //          .valid
		output wire [1:0]  av_st_out_error, //          .error
		input  wire        clk_clk,         //       clk.clk
		input  wire        reset_reset_n    //     reset.reset_n
	);

	wire         cic_ii_0_av_st_out_valid;       // cic_ii_0:out_valid -> avalon_st_adapter:in_0_valid
	wire  [15:0] cic_ii_0_av_st_out_data;        // cic_ii_0:av_st_out_data -> avalon_st_adapter:in_0_data
	wire         cic_ii_0_av_st_out_ready;       // avalon_st_adapter:in_0_ready -> cic_ii_0:out_ready
	wire   [1:0] cic_ii_0_av_st_out_error;       // cic_ii_0:out_error -> avalon_st_adapter:in_0_error
	wire         avalon_st_adapter_out_0_valid;  // avalon_st_adapter:out_0_valid -> fir_compiler_ii_0:ast_sink_valid
	wire  [15:0] avalon_st_adapter_out_0_data;   // avalon_st_adapter:out_0_data -> fir_compiler_ii_0:ast_sink_data
	wire   [1:0] avalon_st_adapter_out_0_error;  // avalon_st_adapter:out_0_error -> fir_compiler_ii_0:ast_sink_error
	wire         rst_controller_reset_out_reset; // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, cic_ii_0:reset_n, fir_compiler_ii_0:reset_n]
	wire  [15:0] cic_ii_0_out_data;              // port fragment

	combined_filter_cic_ii_0 cic_ii_0 (
		.clk       (clk_clk),                         //     clock.clk
		.reset_n   (~rst_controller_reset_out_reset), //     reset.reset_n
		.in_error  (av_st_in_error),                  //  av_st_in.error
		.in_valid  (av_st_in_valid),                  //          .valid
		.in_ready  (av_st_in_ready),                  //          .ready
		.in_data   (av_st_in_data[1:0]),              //          .data
		.out_data  (cic_ii_0_out_data[15:0]),         // av_st_out.data
		.out_error (cic_ii_0_av_st_out_error),        //          .error
		.out_valid (cic_ii_0_av_st_out_valid),        //          .valid
		.out_ready (cic_ii_0_av_st_out_ready),        //          .ready
		.clken     (1'b1)                             // (terminated)
	);

	combined_filter_fir_compiler_ii_0 fir_compiler_ii_0 (
		.clk              (clk_clk),                         //                     clk.clk
		.reset_n          (~rst_controller_reset_out_reset), //                     rst.reset_n
		.ast_sink_data    (avalon_st_adapter_out_0_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (avalon_st_adapter_out_0_valid),   //                        .valid
		.ast_sink_error   (avalon_st_adapter_out_0_error),   //                        .error
		.ast_source_data  (av_st_out_data),                  // avalon_streaming_source.data
		.ast_source_valid (av_st_out_valid),                 //                        .valid
		.ast_source_error (av_st_out_error)                  //                        .error
	);

	combined_filter_avalon_st_adapter #(
		.inBitsPerSymbol (16),
		.inUsePackets    (0),
		.inDataWidth     (16),
		.inChannelWidth  (0),
		.inErrorWidth    (2),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (16),
		.outChannelWidth (0),
		.outErrorWidth   (2),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (0),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk   (clk_clk),                        // in_clk_0.clk
		.in_rst_0_reset (rst_controller_reset_out_reset), // in_rst_0.reset
		.in_0_data      (cic_ii_0_av_st_out_data),        //     in_0.data
		.in_0_valid     (cic_ii_0_av_st_out_valid),       //         .valid
		.in_0_ready     (cic_ii_0_av_st_out_ready),       //         .ready
		.in_0_error     (cic_ii_0_av_st_out_error),       //         .error
		.out_0_data     (avalon_st_adapter_out_0_data),   //    out_0.data
		.out_0_valid    (avalon_st_adapter_out_0_valid),  //         .valid
		.out_0_error    (avalon_st_adapter_out_0_error)   //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	assign cic_ii_0_av_st_out_data = { cic_ii_0_out_data[15:0] };

endmodule
