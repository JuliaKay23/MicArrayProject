// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:16 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V3BLiAk8zu7fO7zdGefvqYVKcpklI6VCysNQYl2KtTpCpilXto5RJZBd8Afdvm94
nV+Lq14mmKrnMfqhKY5j4/XQQZqrjSUDDFHkmtiep4daculsGqLVBZYOpb1F7OV9
6OxTCU27yxyVsdytl8baOClSHoYnRRqXvfTAcuPlqfQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3104)
UftvjxQrVLP5tpz369Ykvq/h6/cT+P9ADxWIa2I/3OiKqKYOrhFwV29kFN/AmNSI
Qxfcz2zm4JmuSPTNY5+hCFLz1td+LZQffBZoNJsXqk4Y4/VRFCRHUicrQCez2aX7
wA1tZuPsLPKRngl9AjhAS1bCVMwhk5wdh1kBQhiYfUW599pajCzBIekMrOaE4Fq3
pxgnsCiPk4XIdO90ufF5eK+Xc9xdY6Mll95NBMhqidPuoZOD548vsDqkpGE47VEj
rsmhd1VA0qFXmmLAJiidRk2gR3j0kFErRCECcLSXmeCrri+bFLWK4qSpmlrb6i+T
Ijo+JmxgoNMbrt5Uit2my03YC1mr6CPJ+h+Zug0kV+5nH2X+kc3eBBuY58pmNsJb
Vqzqm2MU+7HdE0pRSXn4bgqvAtsfYtCqQPyNlrQW+wt7noyGZCeOosXxtdCl6eUb
rQn5I3w5z04NYtcGZaEruLtbRRWHHn3qWke9lk6tfuHMVYy+jNw0opU1RuMyNhSv
/UEY19xeWZdPkPQue25KW7lXXTYLn9KimH1/TE57uyedQEwcW8YvnOm49AyBiGtv
gYLnUOCyQR2aLopmA+QCu9nMRuqJ7sWuxtY9lECSkpBOLcnV8IMcLP7FysD/mKyx
ecxofFEAogQ1dFBGj2vIdqXHoU/QoionU52uP3Y75MP++Z36u/NDnuayCF0T8P93
zvBjS+psadsnCVNCwD6bO+mDRuX6LQvaRMT+a8/66KHWyhDO4bn/p5DhbSXLseSD
03og4ye7p0mbXOUcnDuPTekoq1vJtP+Tm7Pf7yCYPyRgn1FqiDAVfi4mti1rAzL3
fGuZCoS0jrvyawVeKs/Co8inItgIGYvnC0S+8nZh3cw/s/0xyYEqcHqL6jJ50FR+
M57MrxSOlExKyD3D1AyuAcxb2ZVG7M0/hpn2QB8P/Iy3e7EIW5wtdJM51WUtGVC7
fjcSTSug3IYV2DX6RDT05IygXgXiY+6C2B1VEBibKCXDEx2UjdNI78NsBV89njdS
fRxH7SwD0lunTr0ubCJ9gywV5MXCqUuD6szr+I7ERefYTW4FrGooDZEZpo4rt33X
fMKRObuOgJd3OEPZ8tccRXgUjXdnuftRFs3+PXCfOkTGe/c2T7STJcTdIzU7fQFg
F01t4VkkZ1cGnNAk/8OPi6FND0MK3SzcHu+izcxs/kSErBM1tCQI29PrMlPXd7oo
qdV+Db3x4HtolIYmvPlSSuXrWeyjsXQhsIB+pj8JLUGcLRYYhWqhkw9yzTEMXRWH
J74Lq6PQSUSar5cIoLJ2L7+Sxzj++32gQFS14OgkTBpjukHjFp4WjEzJCjn3fEgY
xGBqtJUAn1NeYXMoYTrv1b6NEq5rbGuaMtvHPEyRN02gkgIsEa2U9F2IY90MiH0j
+YJ5MCNN4Q7ME1Oi23JqMH4+nHadUE8a48KqPvHF6QtPpfzXo+466EB36AHBfl+z
+Vv2PbOmwjQXqthKw7Ge2qNi7Mlw3gaK8jyKurape6mcBNSs7u1XSj6t6fVXvduq
8fIQ/3FohJvyw1a+hZnMUs6Fyffzsmc0jn+qpCKx5ZL0PbT6fKUj5NNR2iJbUuzW
NVScMohQg6jIpqxvKaiMuNH5xCYd8p3/9txPwbIRj0haVy/kHr7XKZB9abHinTEs
n9gWR+22aeNIzQgsGegGgBEzUScac8cx2iEGGGtApP8XtoW6ap5XjzM9cWAbobqP
wNLzh7eNI8dL5SVvZx4VJsdhoyOzGurfEFemjuv7zXc8YEpk7pVyuaHhQgLhTgyF
Gv0rHu9n17MXf8DTS4fGH3ZeiNjutgMhS99J/ZgsO2zO3kkWOhrZWxRuO/P8X0EZ
uP7RToWvVEUm92tU+kAakF8SuN4UFVAxBNI3eYRf+a0AAxmY9AyrfQ/2bpnKQLTk
AlQPRxqWbvXFiwN5bcoZrqsBdeOveanG7mv2fY0CKDC01xIsLgH05KeFOHzWYUCX
5tmhJlWJB7QTDUhJj6v2pdwvJ4J7UbxWFTXlG63pO20/xCR/bSF3VIAx4x6wMEcs
NTDs/VgF0tozx+PhQ6UWPgFzZMzO/UVUSk0OD6RoVYV9Oo3IiMsaWmsvAFGSN/4Q
SIG0sOq1m+XKk/7JnmSo5mt5dgbJ2DhsPN7M9S/1VTxK27P1lhiiyxhFui5/Em/n
JtV75CgpXgqVUgYnn436GrfM20aakdYkx/JXwxOopKL1JJiFnZR1CISyRigsg+Ju
rP9TaaLVh67qb41814fAGgMqqa276EBOd+9frCaasxKHXaYT4Pt2UjUI4HjMoDoV
3CRdKNTvRVFPSPTEoMAfoGGj40P8YaB/A1oPXz+pVzRFFLVT0BhDJVbLn2N0zi/2
ZLdicGNlmgy3m9ZlCctqQ6Dvy7bs21QjkZvAKh7MkS7+98qeFDU7HLNqSCmJiZZI
L55OcTyaMGdyG4QJe15ZvCgDO2hyJwW9iyGgL8ZbJN0sXp/hjucC8JNoDcCMWPSR
eCZ6bH3cVu3yntvOxENcM47bpDIDWPcAUbhGX2wY1rDGOIRtk5ndZxBO/U9qLeix
XR4W2Fk7FkiqxKI90F8Pr6Ie6NEzg8zlInQ0iTsBibWMgp1Wv5VkJEbI0dp3NEqU
NIpe45QLF1OtgT5zCKQadEPezapb+G0uIbiOPj+yqNXrXr/vee8T2PE9hLvFcCEw
eotoLktJ8g493pSlG8OERlxkWF+/MCr1mHVlvxbWMN9kjSYQs37tIkURFlaGte9n
W2NnN2iab27NlSiVEKz3myE4CqQmxCK6MdmgMpClhMLVOkRP252g2M1YHDhXdjpd
U0WHLXM2v4etz/QYkhAV1Gljud3bQIoPDjtiTMdopdJSItOdkPboKcA8B34NhSu6
ZC7z849msgU/VZ91d8lz8Tx6jsDwTDXIltkNbcMi4FrYzLP/eCTvvS5Qy5zgUv29
RVHb9WFWh6zpfO3Sgn5gpNPrXKKyxpT0JzdSExHxriuwMMsJb2RhyzXq61PGo0P3
xDTP380/C3vADUipCb85TmuM8fdrdvsQFrtCq7jt1ZttCPDk4w188IWcctAqTQ+I
2BkRMJ8ZNLqMYVjkDgxaHEf7XU8hWPAYPaiNzAkvvwcCaQtKaOsrZMAA5lDhJNXp
8rlkFY92WyMzR0Mth8iZU+w4L9ZHJDKrifTbSCattXC7io9bhb/zpX9BVmp7Kcjo
We5NnhlQD/VP4NbAsktWEhMKs7Tr5aNnJduMOAewcs+b2HdLOZW3jh+vK4xPzDKL
gNfEX+70TYjkJ96pOverfarfKQOqZCa9nNV5dpPavQ/VYAARtlO2y1eCAmMUdwf5
b1slnqf8sQ/QRs5O5msMZ86JOM0E2GPm9AmIukJsKBJh7EYsuGUh6mqAPPH+b+gB
UTbh5ycRRWmC90XRVAQ4+173almRF5XGT61v6sgqnlV3VSeJwPXiC3CX024v/alQ
KGeFkfhrTopJOwszhrAM1IN+456hKqTk6dtgheQItKU3pX3A0uT4LF5A0ZNblfq3
vHxWgJJAtg74nWmrkp+09oar9Ish89UhrUP4Tk+kNbRyDClyuJ9IlkLWkzB82e1V
RtF1u+50uJ1zEgJFRiASdrS1P8jIhIiA+V1B2SJxsRcDuOYmDXJ+2zNsPvSY05Rs
Kum2pxtQdpJYTXzx0rGWw83AZMDyDN3bVVznZVQ+m4lixyiENXd5ySBMRbkGTaqQ
IfkSqWfa7yXVcAE7USjYiETE3Js1une0HvzBWbHKYA1wx8ua/8ucMib+DBN9Xkag
h9Q63Zn+qeVk4GC3D+ZiYezBE1LuNVU+uagjQ04OdMYVN6nqieo/VbXs87tWSHeP
LyrIitCL5VWJeDNCtrZUWyomTL+AFUMpPuMwJQx4U3R9NKNGXc+7ai8LEik9Var6
DRS2D+yzvIN+BP9gWFDWFPZvOw5dAYrOn7UcdvjkDwvVRRGQhW7UPbU+6AZsZ3/2
RVZ7aH2mW5VDosV18KjUgTgmcBWOXDUq3bXr/fRNhdqH5MqESnqUWGnoqLX/ZAGj
prpw5vqOR4nyEKy3uW9JMlDUsovMe4dbmLMKdiZbb/2myv2QSUuSrWCiuQdHlUQQ
Y6Mf5v0wp6ZqV70uaJj1O+B9SduRxYGmbW0WH3cW6kU=
`pragma protect end_protected
