-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HUvo9EGFmmgXc02aXUgQfAGp9UtG9M0O0ZqlQBAiZMVXgLZwhyTBNGpJaL5GWt+22IKXbtEzqi6w
JclyplojDlkANh2yRYvVKUbM2oOciESJc0gCQ14c93eqlbi8OHD+5o0g+FDHYDaWZzpIplf7Bo88
DrPVWGKQz3m4+1rVG/hcHp738NrgMLzIdY0nT3KXW+xkspyPJ0XJ9CSTapZxP78YBuhAe75QZSp3
V0YvIgYlVgGFFGGPeAc/eD1SZGsDf1v6JWhDVDWqzWheR4vUSa8vmVWjjrd44A4LadYEQGYiR2hp
RO2lLscChgnmT2WItKL9PavQ4m9HrXUShARsGA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6672)
`protect data_block
cV+g51AJJHw+hgnkUMHFH3DnDnRqqesNfsTKQ9jDlk86b1WX3nj2OH5hFZd7WPmHSRItczueuFPj
pHscd48ihTkPXu8D/w+zx4KXcZohUF290AJK14yVaFUWtXz7JUInvZlD1yZVRQjoDRDNMaOGrwPg
rAKOTt6Mbli9pxVuNmu7s3ZUluEZqNwHAlTMnRsWCFhE4+TesIIwxxTtbSlc0AzE+7nCX08BSfJj
2qWI697ApOzmQoNoXBagrZVX1EPtbJ4Fpe2NI9iu+FRFlBNXmxFin8EN8SbLOT5ozTlBrVyp30oH
NPaQZj/PmOAXsU9BuJPoJoABUsUOxci/MdzoihOIdd5hoGCrs5Jl2JHq/iKwBGCJga0LJ/IaFUko
NgasFVH10ft504KSpLhaarlRKc7b5zo28W8nwiS3LQOSMkVzYXDhezXC/dQyfVMB6CSKslOn7LNB
wVGOzF+TYRKPyPlmdBLN4PBEnGJvrL9bT7ELiBKPYARKC4ARu79rcDDeONf+x75lSbs1/9YaqKe+
yveAWaiZ1NYRsJn4nsgUOsH4sQ5gc5jkOoL6B90U3R/scpm8yVgNcfidQTuV6xh9Q5ps88ja7Ozy
+Jm2m9hoqYW4/ZtN/bQO0ZxnSPlMbOkSkuNFeKzZinUN//WlHkV0/Bgq9p57iBVzFQZGNvOJwZDv
uY3LqidSF6gu91MNObOJizlooHVpPODIpm9vxIF6G2+b/i/ppvur1etx6dALjSwfIqjcCDZSfQkh
JmuEd5Abe020mWUXP0yBnl939YH/Lc7z4i4/aZY85C0V90Cx7nzy8PLabKZMRm5lDExfggpMPJZd
A4RJXZEWmz2ts75Uz5xUcL/5XGxB1GgRWwiolU+GbVtry3eMt7NJ/nNFjmzaWXFxn+IwmPKLUzjS
1BcjKcbaOMFDWF3yw8LoLUOWkzXEdvLC2evUWo7MscsDj77HiGfl3Zlxq5oWsUFKjjpNVnIk+/tK
4iqa1NT0Qh2OOUt0lt4nMpj8E0RnaNzjeaekIf9VN6FmidOAhx78mXRWiloha5aysZ8ken0QGW1c
PTsSEUe03ctI4WpqDGm4pyXHX5EfhtGqbWxTAGjqG+Q94juM0DYqzHf+ozn9hFVu/kU14nSgQlVR
/XJl0LIHvcbJGkLcBZL0qHh3Gc3K3y3499X23ssAxg61OX2qH3KFNBI4jBKT/NhsG8khKBtQWpqS
QMPTyN35u9BphWh7ptoX3tGdjyCSPSe1v3sqRn2xzjDGs0ZBHdW9/PDLrF7R6Wnyl8bXUn5zDKmY
+QxUjuYFMREov6iboXUAWbMDvmvPXeUQZ4EPBCECgf2YVn3dVu9wektcP7vCmB1FwPOdIcpBLtmH
MTwMjMczmysPt1t/XOj6FZ753VZRI5zATCSoVT+ADtwJjVV4A8QlK8wXcoLrtM/6ks4JSmheeNQP
R7qnz/I33gEnN/pw/9uyh62O2/BWXAnfMY1kKVnPw9yRYHdctN4VTat8ZDZ4R09wvvWu73x/pbZL
c2MOdrqKOw8f76dKmhp0mVkE85e8rFqo1TVRPk5PmfiA9sM73SC20qAtCGvZ6BA2mWpDKEttbY7B
DPmX6TdGfl86uB3RVTyvLGzN+mxBcVF+HycHr+X9FRjNz5U/yKAcOkvPtKayr6RPVVJ6/gH5UViD
YA6j2LOlKu25GDL5o3uKeKgmP3kci3gzQU4rWcdkKJsSBZEliRlmbhQTEYspCsjXD+fBxLzSS7Lo
dizX0ebjAY7b4ImFEn1UDyWoJwOMpCiUBt8QMDuwtlbBISwmju4CZTRa61PlvN/4+hBJ+y8L0OsN
NiOMTwxUFCqU056gAptaRXh1UGswenCZFwhSJ62A15FNvaUB60e0s57qAdCoGNoh7RcqPegLIEob
/Wo9tEf3ebDeoczWk6Flilqvk2sOnxHHt4yaCgCQtefSD9OYXBsU0dJZCgxGBD8WpHTcLEIn0/fr
rN9gEZ6LCVlbdn+BiGu4+knDmxZ0Ju7Rh6AcHLphV2sChrtFywcvqmF9Eqi71TN0fL98NaAm4T96
wzkYfICNf6xiIP2YYOXlCUOK2iNxqOEDj8SVZDy5kJ0CYqoGcIiPQWNm+SDA/b/ruJbWu3Ud88xW
2y0yH6dE2/stgAh6irH3lWhpv4LXl36xk016G4HM4d8lg1mywL8efwWKfmW+TUXp++I/LfFKVUxN
fk5GLizWL/bN7aLrgBgC9m2ScsoQG2Ng17OJNnRRKbMlVf+dmbkh0gX8ce2YesyZsfxhoduJ8RiF
xx1MeKiA/Sgu82UCsis/yc1W7O6eBkGJEZQZ60tHMgffnUCVZPGMYI5EY4KOV6PqD3sSC3eFcWTW
yj0sxiQxGPaszZvqdbFHXGLURkqXMEWELdH/R4xpA+jQYv/+GQ5+kTlw2Zo48jkHAyk/dhM9mqSF
0feev6exnhdbaPMpfxn8StCZmitfkK9Gc9ItSF7ogX3KBAXfXR97ts9+wcNpp7P8fqTEesBEb1my
KgnZHOKAwoaSLf11eBPkaiE6JR8vsq3YmrUzsawQKqcO2FsUlZyBzUSUvfQPq8GJ3sOB1u53xY7Q
g+qAO5qWUDplWFSkLzAN/BsJ0tCO3E5y9x7rvDLPN7mXsAA2NdNdNyD3mhe91vTPRz5UfBuqE4AQ
ha3FBmL4meR1dDKK20KmO74CFK1M8QFi0uVWmD03yIbfPIWwmfLHDGS+0dHmtrj2RINbDxfpx6hf
mEW5/0o3VlAMk5FhNwkVqvzHZilt+dcvUwGuEipZ4Adfe+5B2jf9r+LzzTqjlnh+0j53nmSz+yGE
zJZg10GQVGE/DmCqs391mIqdbGu+UCTOTjvs9AidMNd0l9ngGoiNaxUjG96nFM/75r2pTaSVHum3
ydx5X2NB6xZPAS5S7MQ2dAX+DYN918TYnSblh6glEko8ECWUe+z8nIVwXXtORVtWxFvMxrxbXMjM
IRjg3Y78hdtINFq9RbDAfsaBZaey6fIuZk+s4M8I9WbEC7TFDjik1uI9Y9sD6QoqSqpUfZdN3iLZ
TG+5ds9SgpZ53pumcmvlh5rhzcgdDbfsBwnqXBOW1QTtLEz/bAiAq7o6uN7WzkzjoDH86TmyZVmz
krST+ssA6+NbycI6pWaFdp0P8jpM0BCZGDmMqhOyAK/K9Rcunwc2q2+mrwJ/o+5zkBSya8kE0mMD
p2O1dzaq5cMJ7viUdysREiu8EeQiItbJAiLuqy+oB0tOyL84tiAIrlCBSzk6P8RT6Wz5/bbJmBRe
wkQNV7eZWQ4c9JxvdW+b5IA97EQNnw+u2fz3XFBNDu4HR61Yt7W2SfO8rn6g95CNy5ioALtRqyZI
WHK/8dIxER/OlAIyrNeHpFOEP/nVJcq3g/cVanRLSHMsjdeduk+K+Qx8relwU28e0SCsWtjEToTf
eT09RStVSjWnZaEBlHe3WrWDUcWTQLpsbBiaqic22vE0qInXX1/YjiVzTLuJWapAERCI5UL1jA62
PPAApDdEYplnMAIXz4dRZJAoWrMPQD8eC+Q1ESLkOBTn6TXq5zhvvMbGWVKkJnJ603cTWBjwhvnb
wMgW+6m19NZETMUY5J1ClVxiDVvWiK/TXL09N/crkRhXSiIZW6698pW94MD73NcQ3htN8Q5DHXfa
JMRzesQ2dT1dp4t3Cw8cEIPu5K1hHt9L8PVGuuda039Ja5auzIB0OrwwEAQB6FIYWVY5AumXlNWK
xGOdjgXpDJseM8DOumiXiYbSWxbzcO9SjynTJ4B9NJdiYjwcluGIwg7hP4H5geEqdokVeNzGS1fE
iTg9+imdi7+6g+sn4z2jA3OKNoh71qfkhFYDSLYbB3o+1UFjiFgpAkpUyAUst0V7w1ZNigOeFHxd
s3I/UwCr8ZrgMhFbdA4kfBMu6+yn3IxPjHbB7a77S6SDtQ2P1hjR2iBfKok30aEPQu0eEa9An4UJ
GerpilxPTR0kWXJ2aTrn6exXmRw16FyHCp8atGe8a9PYE7YXLL20vmx5sS/h/r1XjATjuP4tBoX5
lw2Kl+g1YdiiVJ8Bfs/+ZmDqh7rjr+WS5yEl2WsNIXgItZVpCW/2bK34Lw6M+TvK+61zT7Qh0VSW
Ze6KZ+GK08yYG7BWzDvkKsMwMPAdHRk/xdEniHMbpXXkoE6cJ3cJuZjJ9jVCfXvdrnaznXGeioi1
ALf2btFDgVgUhuFuuCW6ezXXaK9uEz3p6ttKc5pzy+qzC8D5Ap7DkfHes6RTK12Pj0aEIpRgZCpT
Z6J511ara2dUhtgxuY/hz3txTkS/LvHcnsRYI1OuKPWcz64FOrcNhE+iNKpvNDSyAlr8aLvDGJV9
5d4dXmKkbrs84qVIsoH4i46WkcaOis/zWCwf3D1B3lVGmX7searGYgOWkGRq8Vk+z9DBHFoohnxd
YRCz8wsqZpL6hCFLbU9ii3QL25taapTO+eJve9EAO7FFentCpQzDVvx0vqrmC0cTRGuAuUu33VCs
gjbkmxGMHjGPxXx16AwctEib1+kcbwImJ0tI294+RhI9D7BY15fktLxyrr1tKLJYwCzGUKux7W7l
fAKsxLcMUM+I+0nejm+YkSbdJ8Bh8u6XPGqoKXQASZFEY8UO6+wWLjfTwyduF5V9v2qU07wHWWqp
NsRvp3g/2HD+x2Av4+F84ZV6Dwg0fGEnVtVchmUATEcjRtvezVFaM/+h/UMxfq0co91kVIlDdAOV
bHfhoCSX3U1P4mFfZS24vDRFALyJXuswHMpVbe8dYbKM+PUSSUFJ0tH8Dv6EBEGpc8nwpECcKwI/
Ijce6EesQnUpW4I1CBSdxweI1aM7yfdQ0RVeobBoYqJnjaNdZFGkIDwBPK/FzBOwdSjOEW+u2fPW
oc/HAmppRm18MsRSzETDhyfwUqzo2JTuBXJOIr0ZqhAe28x2nQnDMh6IVi0Ls0L8wxYCZNeEDc3c
qI96u7kC5Vv4kzN7c8TsyeKm37M3+nZLV8Owe5ttPjxi2ekMWwPUtF9BTBIy2HYKY5126XZdQGtB
WgVGA/2dlrawwwtJPA+UXReMcutDW+L9wGtViAb1uR18jY7DVjvkEFixKH434m8zCKYVqOSPDHko
3WGLJPBrGAmH/DuHI7BlClj3VNW9ejf44HoSiSm2Z3kWkcy5Vl4wB4DrISgj9hjouzZCWoaBdHX6
YlWR9bDTPDgAmggVKqCGEO8zZirRfhfmo6SfRF9Lyy2l65kOK6QZL0q1g8UNAlXi41FFIlEVGtg4
urRV4vO3QD2XB6MkH3xupt1gmgJNowzU6dauXVIyEHsiy0Y6oNjvTWqqA/Yh0SbfEoEUddV5Y5C6
EzbXB+c+YGdJ82CwDjh9MXi6F+BpCS2svrdPJt6MDNrsv8FCoW8QCtCEVZX5/XjADVWWnvdlEHgp
5495sBXZzUqLxpe0PZpEFthfuXlheLTSzb48WflGidduF+JmIbJlwIbh3r7A/idOFHVnLDTycUZC
dYrIq4p8Y/GriFxKdP2J/Ylp5/g0UCTygjirYRjITzxcgiM3u8wgCvblM2W3HDGzJBpyqD+psxjd
SKvoTwblgmf1DJgaZfqn5mzwXq8Fh6SoBSLGcbTXrvby4etPkCxL6oxebl0sTT/6WzE91lIHqp8J
CffFPL1qK7LsF4OdHY6PxWpmVeu4tBZ8TJdbe+po5dkjdt7Dr1dkoJI1myLogJBMOo4mXaXzL9vE
AxYw2yQktiMXy/J64Vfr9GZNJotEiluroEoc7wHW/DpYgohZzBNdHJckEOVwOkCS+EvlyEtgRFnw
ir/1ZaL0gqSZLo4vEAG/mj51Tf7wiG7T3aKUCxcKxMrZe+tjMcHB0M1wy8ACU3yjtYAvxjD1TU2y
31paUy+g2trAz/vU+hFwyg2HbAc+FCcKoGrqLBWgfe9wcMlO/bZs/tRrywB/GvInIi2LmHFk/zCD
pvoTawcCLurKgyl8dL7Oj/hyP2N1I5cKBqcBgpVmg34h92HrBB8ka4MB1wRqsQjXnygzWMAzFXE3
1Ui83iVMbqtWQHKQwfBNJfn0D6j7U1gAjAZSr8xOoXNbbnq52RkPq7duMJQsajB7IHL0aRIDegD5
c4XpGBdjhBOZEVH4jWPuCBEqq+toQl/BK5XnxFXSdrg1cNarqw5Inq2Wvb8LL2niFClAGEXbYUKt
W+j3fpnmYJkCVlzTbZnBKKXFkqS6/c3KoAoMAlDgaFfzGm8KY+JNYDeOvaT41IDPmZ11irSyn3tz
DTp5RwsvzXwdKTjPIfrZ4Zzm6i2ocVrpCk2NL1wgORHzdtzY4I6EhGB1CC4s/hN2xzCpgk9/4jxY
17IgmM39jSja/DPEUyJykCXsUr+Dzh2sXgv5VhXd4Lsjtx14zHEaZVXoUN8bjzuIzaNj3g44ACh9
gjCAkTPxIeyr4UpV2LAJdxkwyb2j3K33PeVFqTXU66IPgIzYx7oaGY9wuyDjq3ZfU3TiwckNkn1v
BhmnJhsKk5/w/wG1+WEXk9mI8O8eR+Rf5FLt0V17fFcj9xuA08t4GohCpY0MEMPOHpUPtMIpjKKu
veCu8WYKbGl8BwrbCYwhTek51jxYGq1dRzn73Q8vbpSt6sUhj1CCKg8cI4nzjMINHHG0LPBF3q0F
enWsd7/CLhifeneuFclvHgQ6MQt1mxjNjrfywYBOjSFTXoUtHz1UvfeZ8weUUDNv4umdNai3JGF+
UqwTvE+lrJku5gTt05RZDYBCDIrvVrlXW08CS0eCnh19f90Rfa1z3jMFeq+lbJwb+fEaEnCJxOmM
BueRLtKX2rbGY/N8xxtkl8q/CZmuzF0DmmEKztjgBGvaiMWpMiV/LwBmp3LIG4e4LTFKG7mbdjtT
dzdIQMJirF6lajP1zD+eFDToIcJ/vEav251cSP6vP1iM2/RnWW02xrCv9sIzwMd5Be81IkQ+ObYX
5lA8gQDbLedlPM8TZqx+XoiYs2RinGaBQx8BhNNjNOYEXevfbdNwnxR08xplr+rJ99/KZ2hMFw6J
IXRfG7V32+jjmguyTALSydAr4rFcG+ncrnKtIzYKMVwYb3tWEkhKCP6NLLESI2OkFuDYsM4Yi04E
glDc0NPNqOSprg03R8qQaEQL+ob0pXb+Y3cD8OpCfc3qDiw6bW6lhoru/+oZ1Nii7DftPXW5IaRe
6srBSu34/6e9qGWV2ZEs8svXg9GldM7QVsPYro8H5VRG/2+loEc7nHvRiz4kLX6MGl5Bciar56kO
iVHNcJN3pwyExShQLFpjQFNslzTt/AXkOIYqh4JycdrTEwUBXpIW3Z89OBpz8115w029xdik5DH7
15G81C2Q4ie5sCFXGB9gME9QKrgJiUbMdo9kywnihCSVWeKgXuup1de3FttCqr/5PaH0JTMuYkZx
HubuID+di21V/U1mEF8uPAaLWoRFiGMDIXnamJZ5+Q0xqJzb0K20iWjKXBGGL/mhi/+/+K8VKoRU
+usokj3RZPbl4/K5+7G9dxieLznM9OjYus1dnHQ1W/TpEycQoZ7BiYl8ZrWQeUh3AQp8vAt6Tv0C
ROaSrxn/KgKLuGEOYXPVRDz8oo3tqIIk9CkjXK3g+4voyFXnPd1Ah0pFqlzdgXugptyc5hwP0sVa
Y/z95Bg50WaD2pYgQlTziHfm3ohIQXAewITmNkQpJWmfHFbZrAJA/LR4UlBS4zRsxa8t3Z9hMIbK
NK+dd2pNyqGFgfuhh3plppl0ubZ7yIQFOc/2Lhc/AtcEfVdgzytE1pmWrAbaCK+WhIuT/f9N6/Yy
wIfdEIZgr/LkZK5V45XbIsivWh9zlYAnP5x//nK/GLUUiWBsVYIZ0eY+3HB4w4HlhexA3rPr7BXy
tCrSgzDnD3IFH32yMT1Gw3WjYWmuS2YsBMIvPI/o+kggHPdPJBEigChZL/2JXziv1QApkNkIHmjy
DUNTR1Isc2Kv7hwoQ1RL9OYriJ+QZHo/5dCwym4FnrmixoMN/ONBmduNPaRJodIonQbbWQy86TGa
GPs4eky1vh/vuGQrKGuHLhYjxHsEv3j/k5DgWwO9pmuyR5AIzhgJFDKo5oh2CXv4NAc2i4mfR6Wy
0D39XVKpWB/Rix9GTGu56HOJjmvUD0imzM0rZr6uoXMZ5iL/p/D2Qk2zZlPr2GKEqjfXTHdOTKLb
I6Ix+Cxj4w/eUJ/6Mml0r4JkECP7l6xMpeGFVcM11LB9KVecri9gvqRWctViY756EMGgGbnxq2ed
JCLou76jSwfr3xKadkBVi2psgVe7zrqJ18i/kDx3BoGueZH6iwYx3RsrtrziT4ayO4SlxvaEX1pG
xMUYaG6o9WxaO+XD5EIQ2EwnHflHBY+ZGP1TTc9nSbws/Y7VjwtK91zctPnqEqRvYUfYK59c3Wzc
vWrO8HZDyXpKEe7pJ+o089+xYEphBr8jmQHVtiWPqi84egAcQsOumLXk5/UyN6xp4/4TL0GBEoYt
AwHSVB3AmB4gJJfy5/Xe/9Cvwc2AQQXb9W3pDaHZ9M9wwkniAcnrKSj+CIvkyGZpWyM5/hnTOnxY
8UrUQ85jZc29LiJX7/r8nhmDp/HAIf7OkueCfB8cQF6YjlC59rWZ8KcPT5Cf4d9nT7e3j6qKjjeq
9NbGhc54rOb/p0KDySi0cXHoMCohQ3CGB3s8BD58Syxhs/F5zaOzMp3xBwQuLwww80SJnDPdm+PX
sunkXrnd25qLM1HGAr82nzMJHPQnBhfyPjB33YPte6/MV0nZg1wTvS+/ao3WcllWFy06vuVlzZV6
b7tdcFQBHbrqxIsOAz+Ih24hwf0oCnOcQfBAWDufKF20q2Tl8f1HXuOV8fCXd9yFZmmDQhYDosHK
ODHl6wF5BTSX6KNwv10TuXfkvdv/nB7HXgTvQ6DEx3Pb09Mh6WlNNjqynqolKjsizKCfqLLYTF2f
9Piy
`protect end_protected
