// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
x23dt3rZy2J4bxAJGTgS5r+xfQ4ZLlcwoq5AGEVdbjo9oZoszbIMKpog8+Cqh1rCFL+0PJbXbwKI
v5yDdldrwBIMPncV1igZUeSVZeUOYO7sEV/4EoiOXGE83obUqEiYRBEpH5hmA4OcIC40/AZoXNE6
IyL9EEC82ouD3tXw2cCDXT2Bcj5650bNWPzCa8Mk/aNG7qOUSBTmIzXg3SGMkBADGtEC06L8jtJ4
tav5hs2hUoZ7UHv9Uu3qINhvqWm8j5rgI8LGzBwANceziFCj280+aCWfZT3ZU6sx2YHG1q2aumyw
K2b7FYs2vTk7hMMYcKOWjwnKzyYZnO52G/akwQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22832)
lrYJnLdp8uASeaeVPSrLvcJ3q0Gl5HQEteKMhb+VRqOKSUGYTgFV2WPu2r+kjj3N3jVZXFkEp5pC
+s9IB4SoIG4XDHJi4Xp+wlBG0mkdoN7x5IRDnwEv6afwiFOR/mZnyPLSdmWjqGTM3jN7Ki8Qvgoj
/JwyvmVPJ7Ibn39rMyfyz/S45buEkKmHTGn3faDHw+aNcucYoLhO3/GLSp2QOJ2tqJ+EuCbQJJsW
GNpFborZvz5AsyUijTMxU8/WduFSnP5F5JedJbyD/KNAWkwdjDI3HPPMmZUI+5oXX78Tmeoi1GbF
ok5ReY7sjOIWHSOl1E1cBNOMlF6byCK8xDyrrcoxsKEKUmuV2vroQ8Djo+EZVeA4RKF1Kr9NDTYf
2FQ9YXBMIlDTJav43rd41vMK59vdo/pZ9EnpoY+M07GigryvcshzRHhPRLM9b7NuIr4BVbku6ynd
xmWCkNKIebMpuQV3K7NRceq7lygu1CUWSZB/IQRXj3Oz3vhyoRJd4mbgFzo57760b4VtV2n0NwBU
zfZN0My6UOlI4QI9/gpNwC1k5d7w9wp6flSjWpcZ3MB42OkhBQNz6YjtnadDY0+hYr+PhNYjqYmb
mHlGOtDivcsEbgdYj0zpWEbPIWYl6yO1/kpbRku4kXvS8/lIurCU6Xu6NAJ17BIr4VKzWLVR+dz2
XXvdI+pBNiHD94M4uzqJdo5Bmt68Z6k631v5jmhrd0L+UNJxVAIPRMXhT4MRC3/JCi84WcOhU/TS
hjOutlTcct1l/WkV6tjLIcFVue17924bscuGlUPoMgnKusAiQw1DAFRW2CADnhhvahDjiJq+X2Ia
DC0P9byowFT+2sVWmIY4tcPYmaHA4OERqHrhRGaeIu2axXRqFL0QdKxv+Cc3JIP0PP70/+3YhQfp
X1ojlFHg5jb3uaHF3GTKro2sPWHnV4GKqUbOFOeaD2H6h38VzM5IdSIrNhPfPlqyh1Aceir61Zi8
ZDKB0AnaPAEIGyaGTaUp4GPHpgy6NIDAWOrZ1TmyE7ZkixBPlVIDk21RADxviVXc4SXKifF2FQ5+
9KhbGDES4EDxjX243WsmboevwOxLbbZRzPRG5uTcPa6pLms35QzYrYPWzNbPpo0W9FUAzkdKs9/u
X2rGSFy4ua8KWtPMs9VtlCmsrgAA3eSYvZla1U8xwdygVgNJvuW/Pely8lHzAJ9OQepEFOqz8Dfz
ZsE/vl52KFhZGs6FFVx8CZHUfQG95BnGfdqPzIS64f6NB7Tt7IptSZIO0cRklcVOIf+NhaaeBvlC
qBhXVcCTFOJ+p/hQuV3ezURhS1/+sYOzzSTXlFPBgq4VxRNDQxu3XT7cgS8M+m6mxhgwWNVyNweN
Gt/zLBK2uCO/8/ZvfmJA5MfEJCox8ttEFnoz7Tof8+efjYhTMsr0nBxiOWlVLVDPtvdmMLDAjJUg
wXPi0Ht0XMe8UgNf7odR5V10scpWobyhm+RY/VbH14p3AaYNEAijwjOZ6MJDoVe9CFsrcM95D34A
jCHzqxrw+ya0OITwIajnhjIAjn+RtcsHrR4FKRKEfjkulwmS/ndv0ZolXL0U2qGAHUHJQuQhkPav
Z/TQCvYkvvOSK+wSOcAbkd65xTZ8As69vZ6j0CfScOU0DMRkBVrGyhDJtHNSZY62EXJo/FP8XvlV
Z5X3ZUQWxeI44UdrvPUYRohIvEuyA/akqKeJlei0xdTChBw3pUh5yGeN9obURVTEUmwWEr+XUucd
QmNJnBPf27eu84rJitiUk2Atx//Mn6bp4arOPzrai7IgAwKUybTxxCePYYISVO1ma01/k0TqrMZl
XIDCVpg9pmQY/5m96DS8+uTA5a2nL06C/TuLVvBud7MFHofjJYKEmrvyZ/Q+I+ZykzdsJ+mmU9/0
9E+zIXhaHyUiA3eGeiLndsRODx9sKrKYhpgt6XYThJcipJ88q6QkT9xmsg12A9B0B0LsXVIwBySB
PnaEjN/+KgJxRIk7kqQT2ivuCnAZ1oD3J8FT9ldHX6a7ZNgmRnBOmnHpyOyboXGJcx17XldmWHLN
stKdRsWjqozktZAjRjpv+8/YplqNB3aEFt00uiHhbrdmAkHQHS5T+lQ7niFy31rxnvkuBBjke7bJ
PnIhzhObof+Jvpb3+Wbkx8Nmar1zBHL6WQapKt1oIQoHmUXRSGKq6wDKuUS8IY8XNC/AyzvqV3hB
8G0yjSq5smv4BbLbnp2sDUIOXh6A7h8DRmREIGBME1MLYIE9aE9ftJ3TF/NN+N2MahUbl/e/bwLj
k+5ubXqzZyoE9FVRaRZOvzX5FePTa3gxVxXeDhBHWfZudyN2VLFP9WdDd44QX57gawIKNZC11uo7
z2uelD7q6JftXBv7XMQrdTn0WSbOYD9jrC/YVQTOGywOAFKg57w4OKGCQsZZGM9GAZli7wNFFzBJ
9amoRqGH8y+u+J95Mjvzgmgg1A6z/59RLRo+B4S2ZMh/Ris6gO+Ds54dO33Pt1/mR8WrtwAMeHI3
lOen7LVtJBzOYoRRrglXPblxtRvFYlbbBst1+ILSR2VohdLBkKbUcXPRyV65rogR0U+gLQfjmhhH
FDzkHRrUll2xriuZ56ji5qL1OPaFyI0lJQMs7zwdxitjgOajvRbHzK94JXSg7Z4hDncLrJWAPfC3
D6mru6uWXA4Hygr/ycxkGnrDNsFM57FEwdlrh2aU93j+AVl5bjrsC5yfCQ2324kQlEFmPgq+XPEE
9vuuKsU5uFn14CEdJyVPGpo81WunAlmLOTwewVGWcUyTcQjITWN/3jAz9C+lhxE+TRNJY9iA1co6
oT2oDVGEYFTS8XC0K8PaXiI1bgFOOYxIt0rrKTdSATQfzhf+KeBLSZetb9c5yrPNWXKBQkOn5/Zo
TbMZexNQH0Iav0EHlHDOmqvFdWdjRryiIFYwaB+UfATbSXI4Wp7hzq1dVvP2oYuZ99QIHnzYCrRd
7O5duALRuX/ZLOu/butNoghG3QINqkxDQLLkcXcRf1Rd4zHwX3E9fCTjS2UmtYJ1sem3v0z+1tGC
d8Lr+XVz98AU10JjaCmHVozF6b36eYY1vgNSGvCx9OSOBCXzALxQ0T2FwiJZi1Zg8ohL2nYFXVgP
c52dehiDIkGRcOAPgNbmoHqu8kDr/1f2bLxup0BITRNA2m3t7TmtXbMU3ImK8Z9xAUWKUhlvcUDL
9y13aZGeBHii26y1aL3bf3IXWXBLG7jHG1Hznvd39RS++S9rloRlqhiFMWQViw4yCHUDbMg61Eo+
UuQ4Bu5Rqx+7er4g3aNSlIu3kpw5z0EDdgiaZGVxrRq7mlzarw7cVoDHS+tvv7iVdkJ0FxEBGx6M
PmoKap9fuHLYAimm5dz9WE5gjx6Po1c3hmMAgN2JB63YVXbts0fj5j2HYHlgZOutpiq+R82OebcT
dN0rvDJHpfjEkHGxXwIe0Lydgim/qzD095Oby1iimlRmRvyVe5ymOb7LUatKorrTrU3MqTMirHLL
WKAAJ3M6c/RqOokNSuofLRPWYE2epw9/fbP+Hu4yAHYynKmKon1XPvtwG2mX3plp4jMzcxJLdBlj
rjM32Hy22evolRW6XSsltMD2cfoW1cwzTZz65Esc28gXm58HpBwlqU7Kma5c37EUDuqT4JcjuYZL
kgKuniaNllShxO5mgrvfI5glablQ30/oAzN3o4pEeFPQH/8D9pxXWO1+vAEdOYdCKLNU6y8JZIxq
xdAePx/sN2c8bjeP6f97GsymysaznbZZ2uazj5ydOVtiUJEn06tZhUde5W1ceelaSWEK6ttlNQd0
lPcqnchb0cxma6Pk7xC0ZTwo/F7N68BHzuaXA+glGm+gVPPBNqUXQJYsDrRbHQZRz0q7z3W6BZi9
OqtiyYuwiNZM5QQcaFRIN1bETgxgc4hS1u0GwgIlj5NqYcTlM/HvxmSkJHacPNWsrDXduf2caLnR
tIGKTdmOOVLKQIPvcHKN6oyTf1yfwCO3spQ7RZcACyX/YcQ8KAp7SyfpqjoBjRgufCSr7ZZPwJjY
fQMLMg6QQ2tKPdZNBBZVP7idMvT2HlgLdNONxX32DHfjYjWpy9QG9YFIVmly/nTkk+EcJGQ/IV3Y
Jb3zeRYz7eiX8aiJJ4S55vy67Wca9fmJ9mIJBiVqOB6j5zP4AFRxK21iHu7qAhbwcHkVt9oV4rKc
ALrzxeLL0NOq3CR5oJdYfJ0cg6DBlGv2d3ASxo+D/Wk5V5ULatwC/g4LxmgpFk7SSi3piy/H1qmQ
P0ZbVl/xiIt1GwK/whbchyoTNR9Tfg4ucjQ03QAZb3CokAFou0CgTYIh0tDFmCY8nKUUOW6oW5FU
IAngKdAnYccHZc3xsQjPrJSQZZzt7SVTpyBzKFB0FWLP6JYg3BdxPm2y5qhX5sKPXB4vyHNwNTHx
tJVHzn3W15ZU40TyIhBs/739AYFwdG1BQKPgoFnH/k0MZEtnPPsjY57YD4ltIrY2YWv/fo7cebOd
38DNMxDNoHxYx7TvUfTbI0E0jEWJAS9r9n/LBsrFKYqgksPDpDbwMHqd/MZa67JXor6w2QYdTWHH
lc6VePp0dH8PMZGAMGzmEzb14zZTqaL6mv2iKTC7khYLxDYLQ1fhS6WTfOqVyVJDbcM+09ZXw072
3OgskyJxiiADpBqPT7qHh0189nyT2nx6a1mzNrnZUs/tvSPRw9fYZoNB1WAxGai26N5BqOHlJIRt
InZW9mAY2E6/6/MQwQf2b1/qDV8nERZtE6Mban9/saBJeKRf9n+OxCVlToRLiGFM9UzofGQXUl3R
KMlCvHooyg47Ttxe9ohzOz/nzv/EwS+9gm7zVjUAK9HzW0+jYRl585LO3sX+pLAy4XGpOPsDT7Lv
E0hajjb9T2VGdSNNXcGmX0WSUDOItyStPBT1jX+NwrjIbzGgxDzC0drKEHnsJLaRDJZCKO4/DGxo
G3qaZVXEPKxHotNQYhqBMG8jFrlJ1duCyjhtC9vjumjN0m4ejd4tIFOIZNE3EaiyOE+yLB+YQKvv
FTw7cV+i/39GWw86YVj9Dy6S9bET+zG2oKN8C9RN7cvT82QV+eyibH+Zqu+c2gY0DpH9JjcVwe12
Mx52FM9oOqUpdzAgjWhjxfRNTTpqrl2wLkP65mEYz1FhYPjNSdhH3UPTC7JePV29TPZmO1pmi7y2
zXW3P8z1Jq1KojpBiVRg6Pd7jdpjBrWePXU56qKDzvqsWB26ddBQoiWhmHo7b1/hYbt1jkn39yt3
VssmgKDqA4hKB8JeeJGag6FuR+6McP093Xt1BWBeyg/kIW2fVFv33ZIWuXdTuwNIvYlhzBz8TRpy
Uxd9m1yhvHNOyZsDAU4hOdMsSi6+OR7I/R98t0IwGCYwnntvGVg82ImwqzO9BSYvIKRWfkEDE+Nh
gEQnwF+hiXxSdQ662MN6jOHTC6SGbDJ1h6g6FyGK2vXrYe0F8wUNvpdlWRkMA46zzCB0vPKysFB4
dMsnERYsPPCrO1/SYC7kVftQMSQMQBg01F1bavtyv1KYl5xxvjWI+W7yMCwLWMSIbtx8kTA+3E9m
nCC4ZERsy9kZhAK5+ndTm51usNASGOlF0W/oPpzjUP30h8O08T1azxcVIeh/Sk2AKHaoAgKJIeYL
fF65kYRqR4+G4KajiBOELHHKgSkig71dIkUDGMDnwfz4YSBeZUfOnUEokRbp++TRBOpdgw8o5sJg
UgQP9Uyr3tgnY5NcL/C6Y/VBzoyapNhEgcFBPYYkCHAv6bdYiW2HxWc+NObhDOmg7lat3wqrf4gG
fQu+ndvSQN3MxQxZq2xTdmzU1/kNkr2hYG8K1dJFvXIZELNhjGZhBlYLt2yXYAcfdSfZmxJMY9Ww
HsBASP2zK23x1JPZ6okZQA9tUgb7A7B1ihA9q89Uh0aZBt4ecosfqDVXMgan3ZR1TNeaa54iFn8w
fUG7mZRvRukUakosYuIOyo9tXqvYIlz1ytQGYKkRDjNd3pYrFSrbo5kTjwjv0cwTgvHf97EgV1eS
uV5ofc0AdrdH54l/NJogx9L0hi6V4UBVjfQreBgdIa33TDP0FNeRT8SNzys3SUWU5u/f1Zm4d+ta
+O8pPOS6JNDJWj6F4bqWNxkb/6uI3tf6DepQ2OA7Z00mnxeWj9k5R6l/KL1pc0MpQlEN925MFzTw
6FbmzuLW8BRN0HPRZyJh2tSEwG09j0C4TyjajaHlaTAGQtM1Pu5sxxKjdr/CaZ6jfzgV0+mccZHy
kdMXlYzu20MiaQRXQuPXmoIVa+0bB2LcE8VjEHpd5uSYdFd336NUGJpInosVT41IkvT+OjkbzYiU
eAIIW9OSeRM+CPlnQfgQYu5OtfYiNrUS3raJWUjaiFaRgIqcJxHbp5I6ENGNaS7gSEZJdtq7LxgA
Lf6I2e0U4UzXigiDDdz/Af+8RYcQ+9adIRmHNrYCtUwPX02iXW3+cUiBL8yssqkITVtBWoCWrJ20
/rAaO+3MWTg0lmXVFQoER0oZrH1hmNAziqq7h2Lenr10YEo8cEExAHjbj//Qz8CR9pBzybotUJ0o
NVRBE9dhAUmQIw0WHM6YT2qBMCmvX7s0g56SwbH9PiRgIzeubssbUD9ZbLLahNJb28GqthGlvgEv
TSpar/BdiyHz57hkDoFN3L/YRzU8XIwZH4rlN3vGyfAro0pSwFWRExZtRKpPqNJprXWgIPF47YCU
wYcynKdGJCQMWjPksXsXQMeBlHBc65ZgB/7gq6+Vama1WktANMwIKTx3xjF0TdC58/1sMO+FEWjE
8lMehjAxtgnXQL4QFPl6x5bF1eejEuNTRNpAZpsF3dN69n8/str3wLRY3RnLra3zWl/RkgcY+D0n
mQu2Siuch+pj5TpUmjxjkOsI9jfRfJvX8k8HpS+iB4irJdj4+8P1OivZMCurecXXSKJEZtszXJ7L
CxqEb8SOEg1/FlEniHazbBeBXKCGB9wNWlHUJ4V/0RK97AIIRcKUNT2WU0hs1wbZsgQIsISP/tib
grKWtp9SPcbgRQNiKnjilI0j3TEDuGPCr1pS56pWozjL6/1zhglk+wForqBfOsOEnmIow2GPfIUR
TJnukezc2oya8q6CJaGP4eHZelvrdX3sFLineYeIeUJ7kLwDYf0k1AY7gK99A0cRoWfgQxpm9DZe
+Odx6DnblKgqJBcnnwE/FfzNxQjVFRDw8SAaeRnnAr7le2ZmxoZMLo4Do3q2t8QAxweyCBkl548Z
LOAHNeeLuTPGhTk8bZSyuulZTmvInPWeThq/Asso8nd1suemqm6+7PXvkENKW2pMH6Z5p85L+PeS
YylTv6MrsS7hkz2xhrWl/S4cEwyJpnGSPU2Zk7vx2IVsGXaeKVz7vqsY96wrwrVMkxqEI3Fv4j2x
Ixpg0atE15WsAUe5/cu23IYs+zMEp6NTROn4VIe3q7hE1FaUZ4bsW7dl4gBkNGR5CPHqmGlKgelT
L4+jfe5ke11VKpmQ855bZiJC/eql3g8T4gC+ka9r6qD/4GBUWcIOmjRXkZ8W5FB+pr7tyyic7GuI
QjYchlCbz5gG/nHHAuF1dSpK3NmhNtvZuajpRZ6+68ie9I5EUdGGyh0dWt7pco5m4lspYMs1yaj2
gFBmaErKFFsoz/LuDBSkSal2k0mrvZHY/WC0zSAqab/yyIArJXIkZCVo9zHI5g383d7OdVncsA+q
d+RmDyU/3dG90cb0DA9DLZH3Tay0RCidWNXvpOu2Ry36EFnMV+wC/NWqnJGIOdqRp7mWxT82x2GC
p1MpElHEmrWFDiy3DuAwM8qVtTYG/loTT/9XXK3Q3g14Mx/H425Sc74U6qCvMkKtQA9acw1VM90/
xDfx1ONcS6WeATVfKCTGcoaN+lmSWSmD+cbMfKiGM9mh/Qd7QVuie3vZ2ZATTNwas8MrBehioglE
LfnaE4P4QI9Zew0nmMgQiWrHAI13WDbiXFmn57dWrbZKVdtV5umAXQ2ww990mVHBBFkb4i/yW9gA
WxUJZlojIJ6uVIyIsGukMO+tfVGzWCK23y+RjjI2ouoNxah4kCLFiMmpPhXBEafHQ3++2a/Kqsei
Vt0W1lm/vyJcWAMPPLqsG0UHMME6YfPIQ9KoiDM2SmIHcfxgOlp0AMR9ftyVlTmIZ5bksbJruLMR
yFpka8eGwejLwc4k6IGAIiRoBmBi6rdm4i3ak05yiDtHI/3Vba5QH7A6N7zGY38Zq0gpivM2KVu2
IvKlX89uFaRHMoCpXkkem5fJXhD6NjIO7T0K/Hv1uRwIaRJuFaPV13avmHQK8qfL24GaAvVCYFTG
FjaerPGwRYkHUNuD552AZ5mKCBWEpcS5sIRfP0pENp0OWKD/sx+gDl6ySIerRaCj2jyDJt4XdlPZ
tAKjYrDHhP0TvSsCAT78DFxi6HDPlT2L0vl7sYL2nuNTFn7ZPUm/Bla62jcctBb3KXlFXb5fFJmz
PrzYfu06dBMAG6la9VJdHnpQ/IbBhGn1LdJFMVA7cigcGO11QrnCpV0icXRO0LkA09TEQXn9YweI
7Xkh6WVWtSSFRuNozyCzYEeGWOMNNW/znCSPkAuubaUcLLGXLJOIZ2wf/GOvEejrDgYcSNS+pMUE
9hAE+VottYj2bl+BQqd+DVSM8TEvjr5k96KoK0TAmgA5p0aeJl7QFI9R8chQ5QvBfPSqqwYJ4HbN
CgwnvddM5ic9+7aBY/9Slij+vKidpFh4IV+5RWtNv0PSh25DtcjhuWFo5nFjO0GupEPL+taNnbO9
2rPsoJGsrNfBvLwaK+LQfBlrlE+3bLuSaYBhXQMQd/YIkr9Gr0R7GwcbC4oaMcXu/Ahi+fD8PyYX
vbFix5oPObjzGXI/pE5Wd3DgKU/9sN2hsA56zWyfdMXAq1s5QOuDw3RZEoeV17CQz7dvhp0nnvvv
6MIb1Bxuq8B5Gzdr7oyfFJqCexaUp1DuNoUGAoQErZ5XsjgaM8x+H9+u1smK+fywBerTIGn+258Q
VXqB0MWjFvSrFs7W2wrC/yTH2lmwiMuyTvFhfQhiP27Qi3woi2yZ8vCM+rzRB3pj41K6Mt2KyjXX
wLOD8vKf8x/D64VLHebDtBRXA1crFqZ8XxzAE///HncbL2YJfA1ZPOsAblQIWDisg6Vj7Gh73Iwm
kcxUEYsGeMaHcVwEasyfzsHEkclAqC5yKzoaQby8hmds41mBrMpV6GFGfBVut/XzQ45Dsbl+wXl1
xISCx7a3ePXT/YGqsmsdxcNz5dGfESdQboSjTqN63abmMQmrTrB6Z8u0J+QtOizMtcwXobT47dAJ
CSd+YmxjTe7ZlQpZHmfH3GMWMTs29buzObyjk9EUrt5N3XVyolbB/gfInHgeiHZI1rZW73I3hN98
Gm91WMQeZRKSzWSe0NMF0kRNGleQnzSw8uke3yTbdOEvkBUkVGIo+yCm5Hu95nN0GJewDmBJffgg
fLx+bTEWhpZEZbRZ9O+kvN/m5KQxX4nEjIvUR3mNQwAA1XHDE7cGZf4IYp5HqGTVznp0uXQdGAbA
yzCaw4on3KrDlxZTfajozT+ATElFr0PAxOC5pEqmWUTgE4YlnESk8RuIKSfl6ODpby0P8r81QVfj
dGHR+2YLdFzlmSruq0vvCCdmY0Kk+Um3H3AEw9rzUVCs+g/kzZbcRRBljE0lJlkK4D/2LGJTIDqA
1MpJwOr2JpFLYjlKOK4i/r7CupY1Uah1dabpVdGchnPe2EoZyRQHcfqcFzNDfxTadPlNKJI2CcPh
2MY4/6eD294fDowBQEkJ3JIeRDQRZrjUjMDac+0SreN6rEBO05aidVzavBRLsHfsO67MUdsBXwqV
0F+gk1WPJuSfjk5LL3FAaWmam7cD3Z4VwnyKOpgpz6Aha3AuEErjBdpPgTZFGJPO0MwW2yFidTXN
t2lEUm42hBVuO0rj7tYit7dTHK5clMTj6yBX1z09qqR+VwepkYKDx0RPF7rK0ePauQEY3Z2t0Vww
NUau240dFyHcj/N5aR88jp4JnZ286gJvhWULGrWZHa28zCj9TQmpXlKPEuROToA4Iz+Ly4ymy1Rr
mu4tY1QOUx/W6Amyn+36KArjRJ77mab7baaeTh/dn6X30I4vigWjZ49aXeWOkLNU7OaxkodtdBbU
f5aDTuRWuxCSTDpGUBB4g7e1XMCINxCwvAzhRkxuf7K7mNO5kdjVBvOknZKB9aMSY9Z62cXrnL+u
DPlsdUIHt3rLVvLL8tdpIcD6AbDdkcOcHS7Z8WGqlalVLTiJAtv0Mn9Wxmbf5l8nF1iYeBu6jpJ/
TrQpy29TFPfK+NZCe2jg3mT6SpaL/Lju+RyeKiIXTQyZFMoxujJkwtFituPCWviiz4zkObLKI0yj
Fys0PZkN40tLdHZGcJN7/nHGnJPvxEe7F5NapHeLkwS5JbAaYygfUjrT+9LllS9T3B+hyG3vyS6e
bdYKRB9sgy8hSreSxuUKONGOX4AOMSNZrzgKEqJAAmQI8DMcNndi7BXNbVzRVQYzB4XLfvtvLBaW
wmvSs+BTFlKq2Gd6/zlxIRrr6lLpf6mfcUh8EyPAoRro2XqkTVXdWzcjuNBhYk9Va8BxhUSKBeTc
Hw/kbBJGSc30jpa+P2wMmDPJPiVYOCzFpBEs5s7qEd6AJQL432Vb5oXCjjSn3UoYrfja2LoByo6u
i/Z83Qv9D+ycK7Mo8oc+Dwgn+plfbBCF56VkGgBho6Ix8JmslxBbQHCZ1no7MmacfiIvs65MI5LK
Qyz0zFgXHj6hAdS9C405dHymFke9F6pz9eT+vh869zI1NJLn84SrBvRc1ouIv9J2YZmpfSU9ez63
ugVgQYa2dVGLHXIuvtQYtrAoSRR6C0Y0qLBLgVsbWrQ6nzhK5y/Uvu+0eE0kbkZ93xfVREULu25/
8lStdyVluqCr1ET5SFNvqBWcE9SSP71Djc+B7b3K5aGGmsi1AXDzYDFCIDngIexyt2K18wYSKNIj
+FklszsfOAKDqPq9RyNEGz1UiJv8owQgsYsMG4n14jBhOnRPgazMXUJ95ueC8KvXx7hYIb4CS5cs
Mf2rRqn/1EAVUSfC6Zb5EOexGFB6OqXQ2Ty7+XEWOLLG6G/Gs66nNqzk5vNZv+d2aSjNQgoLtx6u
1gwb73n1KXsfLnM+NgpzYokREZR04PVfhtGCxX50bd1QlgQoBllV7flJ5hqnqMaWyzhtWYx4JA0x
mAdUyvXSwP/Bd87RfHv0s10JRbSAsDI9myHkkyP9Cbn3HlwnXSSkvffGadm4llZBPC4WFU37Xfid
wvZq2lR0gmIfjhhe/mfLKF/a3CCl5xlq6ImNwHxT91lpuGPwlF2wB9x8FG13HtO1n+gXkpSWPEou
oVdzvfnAs0VwfiTnwOA4/qZ84Beuyg4xVTZ/EwxRGfd7f9qygC5ueeFUEW7a+8SnKl5I2WUVklQp
1M1rGks9M7qTXr+4+jDnlm+QR8chUS8RFR4WTvODdSNoIYBQ5x6eDhQDCcYni+UX3zQf/ykPo1M4
XvUk/0oNzJBbnQbat2GSP5sAV0YTRAll7mlqhEbLqpc/AiyxhUudctQ7SzwexndA1ko0L+tFVlvs
Gs1urUTyUjSCtIxAls1+CFpyod8QKJ/fss5447Vp9kk/miZXtmED6vKJvTiGijrx/xbPkQkTmwhi
o1OnL7p24QUC2G4+fXyl9nsbEhBU8x63MuehOzmYTuUQftkW7MM9lH8T1vWUsAgbMGp3L8HZAwjY
ng28AU2od7wf22jAHsJAKLODBzwe6Ao5Y5LBYnGiOUw/uqqaY7rXLpErlq+AnzZLU3IehHvDaTm0
x1N0hhE2chx13ZBbWXhoYYzbpfnXC+Q+lV3db/DByDEU5xdHZrAGYTv7O4yz4WqnBeN56lWKFZST
zyG0KRscmeDr+BV0eV9osPqDG/bj3GunjiGG2XARkWV9JM5NTHoBTlblKORyTq9dFbmnd24Gn/Kw
ZQlP94minCoWTfy/qFZcG5jPB+Mp9ucWrdsNrqLrP2Mheigux5Ivz9ub6fs0DQ3T45u/qjZfHQK1
Bix3SzKFPuDbZ5aSEZnL9/9AUePllSHet/lyKQlZzWj3+PNO2kd0wq2UvNpF+pmf5GvwMMzOe1sL
e/AjH8O+meZxZKyBc+SdD0ZdRjfJ0X7+94XgK0gz1drHl9t6vJMLhSCsYdD7wBonGSsJZkVPb5l3
Zed70nIG4fKTkwygb3r4O7F41Za9qp/ryjdkl7T8e9QGGSWDFudzWfALXS5u7vycuRVdi3X3red6
kGvxUAL4j1V5eobn0blT/p5vAg2fm7HEADIJEyMGNEts96gezAlpPoUQ/DBzQcZrbon1EH7E4rYl
+Zgo258eI32h2+vbzyjHbCwMu7UtVbtj/ez6L2jGmjIhWSWO4Da4HT0rIAiFUIyWosIaDY5eH0Ht
1r+Eb5BFY3wNgJoJSTMOMJEKnk18w6VjUTbmZueo0VB+GvOYj+e0g7tQ1Zr5KrFXKI3iXTOtkmVr
4vZ3FyXCmpuLOWyMyqYLDDktLVdAjz+fn9KVftMwpqt4VEuu9y8qcWsBc2wA3KvCtjooK8yC66EJ
qjubLRT0+M96zPvLQRGCuJ4BATuv1CB7O5iql0RyUzhdu9Q71NLfalIYMZiKX7eQKuHYvFYaRXYe
z+xTvLgF4x2tLc4e8fF2eiQtycFtg86ma0ETgjUZChIzAwwq1Yao4vrl2JE825dlUXVxHcRgEFVs
9ssoKoHGSxNMmjZD/3m4OQRtuUHb0t3AUYukmS1BB2Oy+r6/lIxNQIn8LMDH3fvEyGGtvGuV4/p4
4WXB1OWTFMoUSN+lduzc1YlUudviBDc1qWAdNZ2m3WCqj9iS33bcD4G7AM8cu7GSoQtJ1uciaXn1
XJ64EIv+ut+MhPUX3fawGeDesT+npJx2sHSSy8xL1r/6tJPHsgyRrTqB6gl8u0Tggqjjdzueo2Dg
Rk7PLOX0nfhmOvJRxvuSGzryKKgXe4hx865OxSG+MmxD+J0+k2FqpWvoZLaNcOSym0YRGeSK1Csk
PvGwAImAu82swN0DjNWmfuhpDqHN+FtJh0VdKD1mPcbo/Ro7vgn6CupM4y3HZRDbJgttkR3N8CZZ
IFLY7M2Ii1wzbrY6NKO4C5BDblI/PW8H0vtjnkuWaMI6jIYzkTXPDQwILpk9GC15KOrAHcz7NTX/
qRbal5O9jv4DSjkNCxXsNUgjFHAKrqbiiBDAu+LBkqciDC/eXZQ96rafUQM+JdPVNPkXn2ynGkMu
oZGkqwIqDBMqFUwzkS+gXiYQ/X3hoel2vkEPc/AMRziFOiLDRHbWkG68qYylKZLDRsgSgnzpX+iG
BH+3QUusjM6O4wVehrCRkOuIf0b2KkSEPI7FMk2EwMAl+w5LUvubrGhr24VliQydjxankUsosAE6
rRV0/TP5DqJ8zwJI4qduV2pLy9hsDscld79PlF5re6coqZqBUSv1w7ufNdEVWUQgjmXAVUfZw4Wh
EDRENTq8niE343pkYIS3JmasnkQWvmnPquZ46ZABtPT4mWF1TDQf9OMD8pHfISRZiKQgUUNvphgM
UEqxOvWkT9AwBR6W1X1iN64YqHNM65opa/gJI3bZueY0EHDwiuWvW+v1t7HuHPl/enCyY8XDR7bA
HrdbqdzR8EtKISgZJKpsM/w4RO/1tJ0RGIIFEcf3W3l9n26z/La3V7ZVNmyOuYVxNea6WZG9/oI9
LHAR4BJiNqQ8fKXkmfDKigLAEzIexupbnUdF6oKjif9Z9zVyUNiMaj2AalUqVX18Rzkpsosfa0y1
8a7JLPAJXTmB++V8v24bo/6sEYK0Tuq4AboYHL48SFu6kYFcM5WwkYQcFKRXKoN/1J/26q1bFxdg
S6/AGD9OA4NpINM17+rcD+A3f4ZbI7SHAlWA0c038RFQs02BOfpzGOQrjUE/EZHg8zKr/WyPKXF6
vMFSU5Xafl9vxZ/uy/NKDUgRw1yVYN8pZKiJqsOBnMqjW7Ckaao+RW+NdG6ZhqM2q0DYLY0p6R6I
RO4VqIOkUb+z3Rj5kIbD2ctqnpujliDwdSkVq6jlu06OKD5ps51FSyJmSZgp3INodeeL0HQwmW0g
0Bqr7kUz0/JhAUrk3T2obKvGoRoeIBAh7nuU2Lj6+Hb6AptUDo+dHETQ/GY3H64oJcnh3PfeFQir
24iFeIrwE+r9Gg8lZDUovD+tTgEGKSNy9aviGKvbpF6cu98+tGaOOOYLeAQjp5IQWESHryW2XegT
cjUBcFcK8WpZX6hKjC6QposBneiiaEKOgZW1T8aFSPel4+hIWWWhAGyLjIewohuX+LobM5+nuvyZ
pcQxIWREKaI9TG4wVAL5Nfo7qbPFalth5pdhBEeHFr3uZHPw0VDSf/+I101QtyzsXCfA1TAjB86N
4KI62hMMIfPBr1GyDiaVCfaFu03mIBW7mk9ifZvv2reGoeE7N8HjG9qnvRXR/4+8CVAbmz4cMtJY
Zxskw4zoUzILUksNBFvy8ZBwmfwtqpaDfjCGboK+hf6XhdXIRnpMNqBXjA9C6zaq8fPTBD9L6H8c
x0+dZ3lh9zRMcTbE/sKC16M+q1gJqZnPKFUOrvXu64pygLJ48GUQQLRh2OPmAbs+SuQq371Hy6t2
x9yr/y3JUS663HFCTYW42Jvh/yCvduxeLB7617+4boOFvMPvaIy2oIn6LekjGCie9pgY8WvfNlAP
0A6sjuVoo6iZt3iFEmqwVJ/+C14jNZCefdEnx0WmZhuXu2HDo1k9JSPGI/u4oRdP4MKiL72QNux2
1Ep2S8mMf5Qeom3NIqwTJAXuzjzEHLj8v+8isxJeqaXr18cffxasaC74zzfgh1ThWzL58/iobTRr
ZmMn9tCfqZDS5EyzBtOGVj+bKnMT8SFtp/SPJLlLDuyW5u9Xi4XtQqaD71efBVyK4MUXi4Q9rPwQ
1a5IkXX3XPuca9d5TyvsAi/nxKDmJC7A87YpE2PV+9kGdIPJ74yFf7nP7E34pGO2ithCJtdjtVRZ
P+ZcSY55mReDYg3sd2bUNJkbPRR0Aw89vCGPU9rTwIoAOlRLOSnp8ZXXgw6YuPuT4U4+7BR22XFp
TwCAP5cYFuFG1CJSzqN4CBfiG8ROKoVJCusA4I4RPou+BF+JUjk2GQu7Mgjfp0lEM97r78My4WBa
BFFADvrtmtkKCEtq7tmcyWJEgHTmLIMs49gHjP6TYvWQMdBCHY4bmw6eSeD3ezJAzQAix57qYj1Y
IYxrwC4D6flwOVRJoki+WOiKcS8jv771xJHw/VVcq+Gsggk8D3xbCsLtVeyL4mxC+oatLHT8OM1q
9wsWPRNy9ZBM6Ijp6vXGK8Uu+7RX9Ju8/8Aq+PLq0QgPSxOytnA6fwJ8HAK+y5O9GT+U541o1Knm
wy3dhyNWYprG5vUvdqhY6hAr3hlNEZfeowCc7LHD9jtATyQF0yvuC0oUxMw6+KYuE7o43JcrJqSL
/fPSf2vIh/RKRTtKLyf7ORDGS1HCtCcQZ6ici9CgqPGyu4Y5NqkDgARhBiLkw1oTJ6Wpaf3NTnVD
npbC70uiYEJ1jPTPfczH0ZEYw53y1YwjasPAlI+UBn7q+O3pkBuSXmuSu25mghFGyfk5oos8lZbe
LY4VrB9bnsYq3Qyb6w8nRs45EKy6CqNPw2YQjfJ8b3vmfgo9g00U34mGfGplli0f7ijh4AUdFm20
k1PDiHLQoHCJHAj3ro7aBqDxkES8i6nziT9eVwStVpgayaw8DA5oFVjJ3OMJ5kR0Pt2VWjrrl/YC
IDgdPzE9w4rlg9XYGbkkGH3CxDp6aHN58g3w92BltFwkr09zQEPVMiQxUSGClQyin/e5NBdEo6M8
PgtACrm24IvAjcC8hgj14cLQCRPWRdlWqKbT+v/59VH9OUFM45UsaW6irGGmWBY7AW6ymykf72TL
015n0LYWz0WVUoYW0YXiIbmRSP8z55GOpqKvQmfkqwM7cukbIop8tOGkJ4NQyfYjbRkPjT5Vf2c4
PrK3/INrPn1nuhMrR1+z7g+YPEVqSMdGXsTL6nITdAwlHCI3fXQn5VTpb/gtvpp9175WpFg4OnRV
QL9KuBnLQ1mDW3XzfWmhzsLbN7uE5AOL45IQiVOb1JTJLc0kqO3JW4T6l0MProIdBDuKN6zR+RmF
pBJCZqjeCpK//9IeXNxhSurI7MnpC8G600Akn3a9LJfgM4P8al0M8WXOfaIqg/JQeG5QwDLSqIKg
F/gmLkVUYMK6UVs0C/6YwoVezy5Y04WRHaT3lpo1EJvZMOhfIHXbxTQ0WfUQR6oEh6F2ZY2hGjgj
SyOL/hgSxR1bxFQmHZAqjU5vSCSJ/aCQvxT2NYx4ukIotJGudAmb0g7ukSvIiARpMLY3qd0/UMMY
NeBzyK5yP5azrHcLluuDQUa6+/fs597Sm4g2Egfm7V4908A+/Od2GtZ0MOeCiTwO1+fwBrjSS4TX
lUd3hSMgNc/LHGZA5Ug+ja94oKHk/FNYW9G678RDnRC6+Dz7BNwrdlN7LygxfBpeujsei464I8Sk
cX8g/XW/tUJvPCUPlWm+Gw0NJ26bHXRYR/sZSI8M7CLSzZi0cl2B9OKcoyrnqZrIAxjQ06Q+aaJj
ke6u/A6h6nTLVbc1jZX6EZUe8Q6AV/trcFPqwM4iE4wlgCXro6vExr+cTE14JeSslDED1S5IGrdX
kKPtapNbLeURQpHoxpWqwANedt8VSZpWkFPEPBH58hInW3vHZYa4cQTA8kTuad4zDwR3L24tTyBd
5Upjmnq3JXj2ZSgc85XKxuVdYivEu5ImtG3c6BOETdVii/w7Swox2jxCFObDDT03gRNt/r+nOhp/
gGvFUyodQiLBCLuHVA2dDQjTQxMtyB3ql1hVNWN1M5d6wjJXcrFS6WYCGxhI+WYI5sviOzRNVmBU
oiKOIl+y2W7wYMksr0oZUCn8jUXTPBAx3wlr4iu0e/kL1V8BIcDLU5uAJpl1ekVv1KFAIC5NjfBC
maXe8VMC0xIa7kl9dHV6lDgTvFOOBmQANJj1kdnhLs9BatEL0+efygTdb2UdX1Unw70u+YbkgRu7
qnGTSLLdGfbCW/6RHnNpT7pTLNcEkI2zF/sA27JQHJnA8ZovgFfa7Drh7Ddd1sUhCqYg1lalj4oy
84o/klSMG5lx3WmeWk4FwNSdN7nyvuvqGwtNp1t+s30BTJruN5wMV6vAQMqvhyUN4ndlh5xy92N3
NYIPf8ZgdN6jyoe/JcJ/CbNGMl260oPXd/JoEbKw1/3/9+9wQU8DDWPTVoPBRs7j/EqypS+PVrhQ
TVZ6ZsqGWLi2Ynz6/SD5V1tkG/o8Xdl1ywXm3IH2Jp8+zwweJtvuMUU2uWOpzZ4stIlU36iqNbNS
JOJWimHlc8Fa7Bh6FJ9WlwTA2ckkO3JHNOjUkj7AhtxPmiWAK2H9+Xb4H2c+tiIRB5e13ezesT7Z
xVoQj3LTWfLU6Jn7IGsCZvdzfrnbGdwPW8yU04hNAZX57R5C/uXAxSiViy1ZnQud+9T42MNwZXZM
D/rOWDd1q7VriFl8GolNnCCLCLcq0xgctYJ505RsDJRIuKVT5SXAv1RYIzkJiXkUzuVG/LLWZVDX
OhXoBSAsrwszZHThFluzuHImXzYpbe5KL0za65tPXosufw2nbX3x7w7/2TUOOz21I+q5fIqkxGpJ
CcKRfuqNo8DXWGde02B+UjJfnYlXSBh3oC6C+DTzVuuQ7OOd0E3t2294esnCTT83azThJaLGZJzH
Ofc0pA5e+FuYHb7PslMTC4azyce7iXf5Tr/DJx+v++YSx9eyPMF4Ip6FyWw7sZO1qUra10Q8Vki8
ele8YIPOzlvaUw0mSSEKMbl45let41KoMu77GdV2+E+PMwLz/BxgU6IwaeywrLFyt7Oj33KkfcDU
1FJibq3JiFId2ShFHizKvnadxuEPMvl73aEul9cl7lOWm9pNH/Wljng3EF6+02T/RkRlc9E13Xa/
Gvtmvy/WtxdvP15D1a3bNnISMK8rW6Q+Q7LUdpsZXM4Ty9su3MguFC23w0DFvcOXe7llxbGfLqMr
U/zGELSUCQjfeT71PsLrjSJywHPnVVNgwL6CHjudQzgk6QyIQcfeMFnM/ivXt75TVmPjLxb2Pn2U
C/tSZhkolfsSvZT5T0YNOK2m+Ao3kHBmQyqN7Ts9idjV9yAGpTLLLDFIRJDn1yFe+xnFeqYIUNP2
RxhWDlAQfZAMfXQ/Q4gIDcBqUQG6KZfuUrp6X5Tat2wx+D+y0CFQK72GwP1q2hRnTHDeAWJKUjgi
4DZr4gFBRAWpqzMTyRgtaXyXTEUIZ1/Ef5dVYHOzsxc2USlYnS7EL85vEZPAVzrVAKlVzkOc7Bjq
X35gFGhHEOvlYoP+mjiZRh07UiOOUUP7xzWrZZSOXF0cskxq9+vT1OTs7uYsoNpa+0A90dIsTEfD
TOmqZmi5svdAZfW6CxO8qVOy0GVKNvaPr41sRek1S6X5uvvpgcwFJFKdasiE0oUDwwPDYVYk78TW
EjIXwYZObAxWXcUb53dl4/QcNjf3Ctu3fbagR+7qK7tVw8mAtmLiLOyDA6Xlpuq3K661ClDcJ1fZ
NWkOsP2KOl+25dyZh0MjyttWm/e+dzK1rRb6MBuQMmUSgE5LjjjR0/SJXWCAPjfcefE+ltkAdvCB
Uyt06uHLaFhiMcEWkqaUHHYl10t3KAF32ygqEfLh8VR5w4dENxXJaslaOJGc/RvX8Bn4+KfqfqPU
j5nQ++9vjMm3j5zVy/sfkfTPp3QOZSESDW+6Qo7869Sn/kTNSxguVSTqT/xXz+0NZyXnZYR8CA3q
5khEYXs41qDiU61ZZbce9/1ubicAVESbf6J7IR7/nJG9CD3yPaTN44mBueqn4olw9ERoxTK8EAto
00eqA7Dp6MO5MOhZM+NHLPkLeibUkGa2Kc/CN8rpvrPaUibn1EpQxqpdZ7J07fmEck3Q7fTaP1f7
3u6KBr9gCpHeB5/jTM1cf/osvpith6ba/ga7CZlJhCcZOL2JTQ3vT5MwBc/C8imVCxFZgA1Bd932
4nEQIlH9CP87K2x0wUmsnxUepGHfwyENQ4g11s0WHK5kaIQwG6HuG0AUyGnVwdHejXjowZ5OK0fc
NljqRKZrOrVClL2eTG7ZGvrSyPz4IWxrYotwSuz4HgR8f1b+CC47J4SRTe8SMzfK8f92LR+bX2AI
O4sZD01/0XE29AISlDs4MBo2npFDy6//RfMc9pj6Y2bXh9pDDJlI6wyg8cXMAuIyIYKhcQcW3zKh
Me0X3tkE2E1HNWP4Aw5A5aKD9aclfR/Z3qKppwT/5HEcHb9MxAv8PNTK5hiMu6ahq/ft7bCWVSWW
Xnihk33YM0GKfJIwI00SQC/h5YOEn8T58QGlC2QMfPw9y0lQFF9/58ydAW80rNTCao70NBHaM97f
jcJ5YHVjXPrr7h75Z3FOmNYwOSLLe0O44dMQ96UBmwN+5i26MIVIPQcuyOk1FajfmVSQ9qIdqeK0
eiKXegJ4rP4YRiTHByxcuD3A/OboRN2Xm+ezmYPvofyb1m9QCUrVt+NfqOEz+9T1AOlmjgycs/aA
iLyjQElDsQH/mAxjttjfYfmXuEm1Sfp45E7VVVr9JFVn1BoZr4ts2OPkxeDGWoLkGOHn3kK3Vg+2
eY/k5xrNcdY8P9sLNv4q7Mj67WJIM1togt/cCc2v4zsoU3PNt0pzjSotFVeq49zdeeHX65FXf32p
YE1OAoNUdbAalY6S6JUldcfjQ+iv9q6bW/Ouc9YjacrLFtCCwRw+I0jGTSiYfs4owFon/8fxPuNU
9tv5hs0iMbO+z21HmHyRDY9EZY0poyxCt0Nm2pCvNm2CJ5TLV6R+wy8vzq7d0gYCsdd9fSGNH7Ki
yEeKc90/fjKNnYq24zLC/0lN4+ra/+Lq9K+he8lSha7px2J9oa8psoTAn214BBm8p+PZ9gomIq3y
tjTJ/BIuNd9nuJzRg5FIygPeBqCVUZHWXWhyI9KJ5qZRUQL0jGGMl54QJN8sZ52gZ3Bs+WAHbC7C
6BplldJynCeITm2w1H02q5SZlWZFsNp6Tm1vMrSUUfyfUVjjpXhl8gTMVznytjiZ3lWpflFm3rJe
X7oyo34A6AxJlajzuyCFApfVbkmNZZqTnd+jvUqKkDfjW0RBNkv7tyWtr52wsPzABHpVftVRfD6x
wyON01obSV5+qTcH93M/tIV8M/LIZwkj1zBHzoUtgMW7/JwmB6pshoBXk/ztXvJspNG89k7pDKRl
ApSxzD3zj6Tg2WE45wFRteZozLJddVx5+Dg0qOOefq1KgI91CxL8blQO/VUYZd5sNM5QuElpsbVI
7wyzCCAwBiRt4EH72mXOaCOPt6lJcv+/LaoSSvPiQ/HPOkBAyx+tkwfpzNRylYPBx1EYXY8F3hPc
SZhbvYPemHw+2tKopARq4g/kL5ZbZUm/M7CSYQLijYL3yRWFvcqOed47nmhRHstEJyhLv/xv1g2y
kky+iDwVOPIUrbBhAxCaCbfA5+X4/gmu7eKCc0mHUpZ+ISS7DkHkzfOsq6g6OJyGJ56CDoavnUtp
hWpHNjGTYJSS6p/L78ZZcuJIUVvgMAtTEkLkVa0Y0wXJCxl77d71NUniHQk9L0HyCs2XJ5/j8Sba
0CIb1v91a02H9jb0A6PeR6xzOMMQUnLpuUakT/4WTOBpXaFbFFkGCvS46cWYZrrTWApKjGo72q41
HzJxgcFUxHNdmeBU/GqRYnjOEfxDEfYaNGTNq+MxCMqIKF6jcqE9/hupDSU5ZdeGtCCoSL4DQ0pW
z52RXFrzd7WklwUk9YkUAPBlrko7vLNIkc4GhiLzjWF7hjheCymL49PYW87ChJm9dX5hCL5V+/0L
nShc8Pv+7KDdYqkeFgXHBQ4xjVrZ+djBHkfFBXJSqdhDIxiMkS2AEjVCN/U24eryBwXlzWRqaXFy
L+sd3joB3jWLcX5i0sdMuEHgtJzG8Sxm31EbLBLGT09LpHZ4mkul3YSYlY6bffqnLBym+F0ut5dx
Vlc3VAa8JWH3qGXWZ6mMqnq1BWDmI8+oxPdz6BMkq8hw+ezUtAgdRB380zDYAGHnXPvHPFh8Teov
Ab1gQoWW7ZWTDmX3EQHF88BCIx/05CoaaHSUv3Ip8Qmebs9MIyiUvTIsLF4yx0d84aDpwAseqnVS
IVIrbnvp9QCpLExzs6qsKz932/z8Y2d4C6ztnKOMG4CoGGc9L1TdzyMCw3byIV9SDxHk8P8qhvOe
RHEKR57Pn+7OyBaQhAcnSpdDbrOEdFh7BRZ1HKhbaO2Py7vM+R2qPqV73nrAxlU1/wyscCHNhuy8
W+efzXW2Mi6s4o8ADp+/+8A2DumkyW8xp8BE5i0XVxKVFhY6vBsW3H2Rx8mKsdNl1/PoUrztsuPe
JXOg5IAIQdVliWA686t2+3+VsP74z3yXOShc3PkbO9KBOrlntvSIfG4snRvhpaCy/o5/YLhNVqFs
Jt8HWGe//t4/R8OXgdvZ3YSBj7AV9Z1REBJZ3u6gpVjELuKwlAzMCrdEwvuCh2PnNOUjXU2c/NI5
0cCQNqVFS+ADfgqIu4w40ffd8xWNIeAaRGcJNH9NlfWpqy4Bjb0R4Wj4Xyp6VjgLyPzSXR1/t2O7
emOS6W4BE866jeJ1a30e8t1bcBw5bnBGEQ+BKMfk/jlu+tp4XzB9fGixnCmwEjN6dt8xXdGnbdn/
r1Rq/D80ZiRYGma088ewj2IoYfgM7FHkiSsV58ZJHZT0RWgpjTKQGuFbNGJa2QEl4iKhL94wI0KH
j7uZZKTj9N7pVPCB56pXRyASRrUVqR6BJeDPu2qJ9TrRaKyUzW4LAAzdRirnnAFVs/4ibz8lbrVW
vP0wO/u/xhAFnS1V42+N3XA4rlh89fKVRwPQaOw27BU9eVc92RiHRwnYyFN7OF8eloD8I+f83j8c
CLdMi2EDLmzDRhtGSYb7/3blbdUal8f0dL2/zaHGxoYrHpjDq8ehUR6Pqfb50nItZPpAdJbBrXRW
DAI1oG3+8X1e+2uQHrs97Dl0CBg800j3ZoxR266W2p2rLgcAYsjwVVdwd7DQ7G3d8iWtqOq4yMXt
QsCJqD5tIqetM+vds7dMGa66O9hMqAu5qoUkqtxPrZ4xddriOgLSuOmrDQuqeTu29JST6G291vTu
npXfeTgSGSxl/uw5TkQOtIruvdBWTaoamP1gmkJZNIPbUx8BqEWPj7ruUhO02tGMjTu47wfbySrV
fZPC9e6HbmzTcDbisjV4vnol+eqkV5SiqJeI/IoRlC1AuAAPQ9jDNd57ftk8MVulKQsTled209qJ
BEc0wvWctatpeZcZ8TeFh+y4wmIJ3wSDOfKzUt4E2qujs5DXPD1KiZnZ5bxyZg1S5khfIyQc4DTP
HRXr4ONid+HEZ0JqofqVOkkL6m1G1BsQub2he3hTtiI4iL4/wyn4rZv9eOnB8myEs29sCAqyWmKl
k/2SxOFRLzvLrnrWfsXBVikhuh/M46+AwG0JkiQAJ73EuRP2QA7Jv6NDrlaMpMVkMjtxxtplxGzo
WHVb6nubzeKX0RRbw4P4oU0UFh5R0dVlV2KZ6cKLUf6XYDQJ+2/oLUs4NuhZ32HAYnTUCm5B1vRh
YSK0wrCT9JtK5foIPCdcSvDo3000OlzdBLz640mdKmaIA8N9aqQfWBqnT1eSIs/glEoAjnXA2KYt
T6j7J+MSGJWX+1UB8B4rl122Leoh6glB0hoUDyu6gnwBBCJlwRjPOz1X2R9qFT7CBKUxdCyKMx0D
yut/f9kb9f6AQkh+Q8zXI8fjXuYS9GJ2VPjo3IInM5YIE1oZfVnm3Pj22yqdQr8h8gnIFp4Dn1NT
JL7aqhvEBh8gF7ymfuMUe6QLTlKs/CBNLlsORCsqu6O/7JyHT9By6f2n2bYNtWf9jF+IRXzCxRGT
vdJHxz7F0Kq34L+O5aVB3H0u1OV4FpxO0MW83vXfLkft7xwR0PmhQG//cL8ML2vQ0Jlrrob6xJ1r
JKUI+zrr+fyDJjKAufGy5kg2qf0Ieu84v3GEOzw1lrT4siKtjXImT/Aycd1y+GXPTtcDzj2JcCNb
ZS16ZgIYZ3Dg/lNhU8+j01Lpcy8C6AQ0WVCTG2J6BG1t5RdF8M2udDTIdl+Ej3Uxq/9DRo1BkNbY
E3PipZDbCkn7vImo1xMrMSB0NHpn4aBQEH0LNMR6itX2FlLt02mwuAqibNhck8bSwyj4rjG37slb
63KUkRODVCHc5QsLIZ3wUwUE7+bwpF+zAJtjMuzuOxLeLsB5oVuBdqSYjZkFf/bTg96LVpZLbWYl
jCod/OuTsBlOQQDCOZrZ5VhY/XdlwBR3ldG3KWTSqgUuzvdEMmHrLILeOxxMksC8/jyL/C9F4A2N
tjGw2RiXPV8znwiKch2MHPP3OoxU4aBaI/PqB/qSe0jPa+t7wpE0VIQGtiQXeMuYezM//frz24xr
D/ubOansw5Jpg4/BXca1h1vcIa3/wMcN41s2KpoqTrksabHvaVCCTpxkWGUgRYBmiCyGs5vCufSq
1IZ5m6VAn1W7kQ1+hOzRROSAzb5T8l0aVG1EDWAuxuxzATQbnt1Lm/qpQnLbMfnMXpNoaalYAah0
s+EDGIHtnN2UoxabgY/E0WwMDQKdFTAM0F6DNjcSh9uiIO9BS/PupwQuzy7zydjrmzFwJjnyPnFy
N/jyMIf2pwAN1OaQSnRry9envFrcKWqug8aSd1C68Jop9Pbkg6nKIl6K9YIcbGBaGOo3ao8mjZ7x
HUv0KjdIAZ5o5m3RJDBiZ15NviI4O+Zz8GfYsBQnRXJJx/usYA0TI7hTPuP8X4K2MF6P0gTr8Kfo
uL48wlnP0107EtUzVbEdCEjOoBvMJYiy1oNFoGpy/hXN6odHxN3bzUyIXZnhD9HzQTw6FuXNRTA4
r9lD1+uiW1IARrk+xdEWeIWUvosiM8KQTp2XnVKyI29cwYWfBV+O0WWSLVwhGXxFNTZv+dXcPek7
5gKSPSQSFTD02XxCP9EPyS2fW5KP5Dat1uMYen6t9mpzlgm3v8o06jT7UeZIKHvV2N4jp9zFWcWd
wEND+iU7YMKgo5Ka0Ddarq0To+IHGpHJmjhLTeYbxmtlRblvxQEnwZJKJO1XeYscK7hlfZTrbtJt
vT9C0it7nFSH9bZTdjXCkLe4kB4FI2IuXMyFyNlPFfkv5z8Ug/gJ5mGAMcbYi6i6hpsGZzSPAsU4
fScrfocSSiP2pljWEOQfroAH15/4lYNPZDjksVFv0/SmR4MokBgunQv2XQ2eZ3YMVzL3Su6aEHYf
qdXhe6hrBsrY/FbELODGCzG5EQ7Kuf61KhQ7EmrU/UD8aEjYDLQkyS9HvRnuKpHTdcRLBcAG5VS1
sYiGFLrqpKiQJiqOggC9GISFtn8qbxje3AqsQcRwH1b0BZM7jZ4A0w3qyRiM6Sx+pOw30hoMaOMQ
l6HcLG+r2q139e9Wv1X7lSo9ZWPeBY+0fHnjXLswJPFFzunPQ+zR1myVozCJrYUpEbCDgxjuoWYs
UIeL81zEX+gW5eSY3lQKIEm9O17M4Oy6K5b/vi0yl/dgyfwfEg6gJ8JxYIiJca9sZVBselxYjDYe
3heXUeFgzFfgqeakMsNsKwsDj6/RCV2jJsJ0WXDXKq24ogjAA/4p/cKWwkNBH1QE2z2LStOTOW/f
gHuR21eyGpY2oXD1xMPp9AX2m9i2un5E2F8ETc5XgLVPrgtS4ZuMC2pUKlxYi52xxquQFKUQXi+s
ZFWmK1KRYpPnD5l/MdIv7XdKQgxgJgpDrU8imsbbds4tIYOdwNVQ+lEZS5sEAtnJzACqiqzJTEzX
wJ2ZS9twB1LMCjXMEHLaoQM2Lg0TWuovbrgAcRaMpv3QPDraiBWh4t8lgLgfh8PKKWO+RBEe1Xuw
0sJWYGU1pwYpHHhXMxmHHpQQvdqh5ZteK4Ms0cusbWTPSLoBiFfCsRM6nvdpcQcWOJEKCRZlonJS
VssFper5sVueW0ujHklM8gM4pQSGuB1VaafjT3G7p5L2sGDXHaNRew//Jqpgw4qtiO2y1xNgeViS
sLofJCEacj6AQcVO/lDHxHSGk3bi7z2tfn7lRdok1t0u+HGl/uyT8hg8EO7YqlTSLinTTVUATkBt
cSTm0I5Rjy1FPgTnYcNKvSdkmBrTzRHRzK7qr6Ir8LEp125xSxM8JMj0ycQEoZJKLc/6NLsKUcHH
8vo4cCqCfjSIybdsVk2ds4sn6ISd62vRamD8R1Q3qr26nL7Vg2qUAU1XDZtVbkvQiB1jEtYbEtvy
OYisfjLKBBy8/lA3blMU8vFUe+QAcvtz3SRFbm78lzXpPsf8f9WFuNjuy4Y9MB1jEtLYay1L4EyY
icHwlG96B8vg99KONNqyOvhGxz8RjUBNucJcCwbzGJXGFM9JFsyD0Sv/bNz+fz4icb2+tCfVH8Jx
ZMryjoJY2/FWpYdhEZkIceXFn48z669JBwH8W3tr3Osj+X946aVaFaq+kCTlhnlmkvtyOzIp2Q76
q0ubJbWfeJVQraelbuPZO8lVMfwdhvGnFheURDTUmJNkI17jyR2JNXMsCb1WRmLbN6hhokoQZ/6M
sYqvsAjroVU6ZqhPqHtQ1xvUP/2GVMaMuUSrnXtezPckpI5wx3VRjKPZRaU18+JhLRkmBUYcHCT4
6zSK1cjSuPqu6t1DvYf1IvSwxS6YAEZBQ3IArfJuLNZ6sapXLtNl+/WavfUj7K3d5rUDWOpTfwyX
Zj5gtvkQIE5Vg3TUejIouIb5c4oVrfQJUywsn/N634j40R+HjGNJ9nJpP4HtNwe6G0VpmYIVtylk
DfyrF5Y5jjLinkYzThd2TPlxacdISfvdh6OuoOhuEY5ZYGYhISxZiovCmttQSNggcvRtWbMr4nGV
O1v0Nps1GHExf/lxeaOiLFalp/eRZ1Xb9gFzwo66kHAtSb2rWXfqBVyuvs3V5bq03TNTZB6ffNRj
NakCHZRJFHFlN4Dsvz+JC+uj1Q3CR+fsTzDuGJD/AHSVZQJAqNu1hv4Fg+hasQjzIPzPSYlVPSmj
BSRNx3CKjRVkC2+7yvbG3+W3/bP3BW1hBVbya2kIVvLI+maKwXjktswkZsz0+yoR0I01U9bQa8HI
t0SR4wISSv7h5K+eWCd5Mw04tKOBc0A7RaKr5yl4WgvjwDK8H0LkYXIYH8PXZBuEaLyMQgniQ66s
VgAoJmnjst8uGy1oKKoBTTU0b/krAb/tvUtUZRWXTPYSlFY4wiQ0lJ/ejNu+beOnv93xi0ooQyet
0FKmy6aHvhMIZkEjo+dUOAxyIzqfieGAVTtENDeggt+BOU9RaroGlAqr/4wd0LrgqiHuQWEcjZBJ
PcIKfi2jw6lu8jAZc0LtcXSIxXJBpjcVIzujf1pbzbIyLBpAjewi0Oj6YSE54LhpagabvZDXRwma
EE6GslQSY6QHhB5JoLxCmBML5P84WsqiqKBAIrOMyzw24ytt9KFFYpgin9OF+nGToS1z8oIyUwFW
Vxpnw4CKGfDKwy4A74pFd1HggYbbsldSYp1AqTg1ghBEKQ+pT8LKs63UjdJ7bzSHAjQQlQvlt9Qk
keTopI3sdh5AgMQmcqz+C6i48DK+eFJVUOR6U/q99yIQsOxciGTGcQyM7BL3SiAC7/rFYANXvv36
ucbDcnvRU6ZHZvZ/jSyl3GnWyNrVSuOEhB2H7dvM2YnBcRYuno6KAsyKeKojt7YWDPZKiwioyccL
bUQ8NNurEEt9RJGekOpv4EhDMaCBb52oL8X588hlz8oh+npc4SVVGGd64joW+T3/+t1TwZX1Bqqt
g7IaPnvCEstOBq7Qd83pZwRk72mvw0TzQpkesyO3ADu2fBLcAh4uVsiuhsgA3MNlVC0ekHenvXup
6C0NUpI/XT293bZ7iIBB2cN6JIeaOh8vbuIm34Psj1ZWCcbW+1nqMaoCAYEWpGdE6CsF1jTysen1
AaMYh5UtNZd50pZUNb/wTJKaD0qB8xwXxEadLxcAaxuNqYV3SixdACVDvuqjdVXc54517Vz67n/h
nCYO2kRCQSU+uyW27prLOgnlBSrNruvq5B4Xoi3CbuaXEhV5MwQWRnqbms2zKalOzgoKatDJ+FEJ
yLq/+0h0yqARdfwxRsx1m2VQkDBIh7jH06YjbxaTnzLn234z+12/JB8b37A67/945Gk1fEMpZrRh
cmm9yKJZmbmHdFkeZ4irjqcGtREhINhVJE3zghmOiGiyX2Kn79jTRT1xQi9kvfQyJIgl82VMdVpQ
Y9jlR1UtWXpX7nUttYCt/Wc6hxYRsedJJLXZtMGa4VbWvZEa9kMJ6yimhGh/ABK18doEL/ywUoAP
ltKVIx9prxIYl8lN87qXFNZt/ZEoXuYIjF7JeVVR/rqERP59Ao3wqe51FwOBEm/0TrgKgH4h1ywm
QR3yvdFxmnDUPFO1hHsTCBpZnsdu9Qgn6hAh3//W/snJeRoQkqOxA2Mgf5+1sx49xr73sPKAhQSb
xO7WqQFpx/E2mVPi2YK9Drl5DY/Zj9bZQJYSm2lH8zASQYB4Xe+jTDg9UciKHYYGNmvhLAXPI5YT
yr3emaso0FVWtpQkUPCmboUKnBC1S8knpoyxQ85bxTS3cvjOeXLu8DycHk5umDx4TgvQUCWf2r7c
KMrVeXDleBi8IU+SGgaHdBGls0vhImJmCOxhSK7WIucUf2bzzE4ulSonG/w8LoHrhXXYVMoeXJ60
yTp6ldLfSHwlIDPz8ET/m1aRL5jpZI4XjpMCMR37dQo9uKY85XNl1uNg9L7S0pHLtJH5D2JDm9wb
NGiC7T85El2SCG2fhsPXV+sWZ00CiDU9kHr7wcSgcWkSSyCAR5eUNdUgdXGXO5Zp8ujcwK2W419r
pmIv38uJfQVEtwyNG3tV4CDzWJDRnG0PAavjOe2HFMrekRbWv22X5oyB56+iBahsxfqegvfwW6k8
bKTgs05YdLMlycUtPHMnnu2e7WrbqV8j9nzqUYn3uiqqv0DK+d5VqzwLSOANzYcKFOE9E4cf+AF+
zsIF1PrzC1oo2u0e0JCX1dNOXov7JgvEry+UriJd6Dc6DN/xiTRcjyPm05BVDw3MCoILZsKronEW
/L9TovVwMoF7Kp1X7fTSa+3+64JscfZM2YpblL3naMx4HCg38kkqQkzNxK+2/tcgsObuHA4Hviy+
+sUYYEwEuSi2u4VQS2rlt6g3nLFaacap7ieiYcZe0uqLUhf04nYfxb+H0uAXhzp5MfYLQikMreZh
emWlHY+vB6ZmI50ord9h9hVLXC3cMFl2+SHrELKdQP6GWLzgCJHGVKshdMAUdV6bMhLTUt854XiF
6MUHz6iXpH0nXss9QKHBL+JmS14FjbgXusvdChRmCrYq3iAPXjjcSvwb2WQ4N19Vme6tA2ISqJNQ
LSl2Qe/iyoN7UtCNfvdix68tX0jv8E8Q9fZY7VthI/9alDqgXJCBars78kV83WIlpcCuxJhPxu5C
VAWLoZXXDBGj12QIHO6f31EW73GA/7jBIVQjA40SEtEe5LlycfkMsWbWvugKP1Tmnu0KewzORDLg
zGDLzf0XjkBgt2hrvLVd/AhGbUO7H2nrLU43sJFztpMS6XtM6ejX/UzJ1NJUUIRQIsBsfCkoC2BD
9A1OBzgZcS8oK0mOFNuqp9/hj95xJ5SMNrVYVNLR4/9h0Vpp6ypBvGFTxJx3O8zPwtm9WOxcUMMU
rHLVQ9cBfvv/UbRtZuYev6ei9XfJq0En4G2SDjaZUpiBOd84tNXEJcbWpF+6EUawY4+RyQzhzm+I
vb4mR15j2gHAmLC4NVBk+8Umw8bBKTPwIdrno0MDqQOv8b4w8Xfyn+nH5Hc2ZVrA1M7diFNrCDpy
xBqfe3Dvmw0542fFPA0SacfgoANUpGIhYPc5xSBBMPOFtM/wrcY9IwEhzmSRWytF0iFhQjsySVBL
BHT6jKHnCNuz3nqrfYWbLOBIpYIhys3cByBRkehDrfFGx2IzZnxaHkA74eNmZq4XJVaSAFtJ/f40
J6YhYeNtKU//3NhW5t+liHvNPTZ1DWQatMGGJO47KeryM+wpJhAc7vd9/15VNrBXPfmq+333jfLC
HLZu1VTwGGRluWkYfDFcY5gvmV/g7Wx8EhawXFOiQZKpkwipFvL5hPZQFhVxOtmzYkmZDRNOXFzn
3/RP7rVbI6C8lOiYqfa/mvPF0y77aOGulN5ZOJj1vtyQh5P36Q0TT8zqkONtkI4Rzdx3zLzOZvE7
53Xc/+e8Rx9DtlIQI3/LMY/zk6FKpolm/4S6bPwW/SlrimE3beT0HnylytYqku4/hz5vXJSkaCR0
fg3MAH8pvteFZw7wZs+rGMKKcCg1YL2SvYLKBmzNVxQX1OypXzfrM0lFCe2ItdxLVqRLAsMdfqWb
DBJK5Xv2VF62HO8q0m32A+SNbnZ7eEkPfGKOmseStQtdIwUpNGZhv/ntVO9R19H3atrcjImQx44Z
KZCt7AyrrjXnvh+SMtxakWc3e5x9sg1JkC7tBwJsCzgJPAEQTZHGrbg3XuSwVTC5XTlN8icyoWS0
jCv2UPXw8AGiiminJKandxEEFYjdEcx4o33Qartony9U6+V1kCQDT6UC3BZwHvOYaJGnigHVY020
vcTcNgrSrTcVT3CAIznw7QzlKUqexgPjGfrm/VWcHXRtqtz6uv8CCOvRVFO01xclxGDJw/fkCaws
8y8bppOgPg0UdbrLhnMdD/aiK5OcQ/afGA02W8XVcntzGGHi7y/2fkgJvOvzG4dJZ/iqFExo9YZk
IT3O8u2k9cnYWlegZ06IqCTi0niRC1Sa7jKKf9COF+OpgZCH8XIcRrYUkWl2KK9n4yh5keOdEChu
2WOZDk74SxT5Tk6WAeXgwZPghJ99rGB3aHnuFvLEMkU8zXN7byMWQnFxA2UySWz8muqoZwYRNk9B
k/AnmRbC82sK7/S414is9VuSfkKDGK3/SczdRSgR84AK4/3Lw+0IS9BbkmBMpsvWp93Xhbqhuy+P
fgY2We3/eR03eY1Sd0hacvHFBPvgd+A73i3JGFsdv9lUl9v8NkRbIbah6F79/DIzmXQyFET0j3uQ
ZNupuUvP082gSt0XAj6VwGnfzpaGKl+cBm1NKfwvxBU1OoYdmN529FQOeMHT6PQ1Si42LaJtR0xJ
bt4YEji3QveUytlqu60DRW4Z4jmK6cYvRmjZMVQhfZLdZ7UlxpR6Y+xQ7wMtcqolfovctEEG2jG3
uaZND3rvmupnd8+/TRpNJoT8ZD33OwV117MQYDG8bQszUt15xBNYyoKmlvEJqlbo83JvT2WFVzpg
VrF+AStUhyDfPRWIjlhceh949ZMJjeMkqFty/HmYyuzWfJUNCbrmqsxCaSWjOXGO3DEiw/XIjf7f
A1TrLlg2kvOH87ye4OULuJCGuIGlRGFBnB1fszbi9RSMD8oHf4FTMiZtRUOHYiNoaXc7I3FgO8Bx
S/tlLVmT7lV6hydEvCxcrISdEcBamBMsVer1RTsdVgE=
`pragma protect end_protected
