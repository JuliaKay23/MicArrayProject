// The top module of the project. This version is for simulation and uses
// button_debouncer_sim instead of button_debouncer.
module mic_array_top_sim #(parameter mic_n = 2)( // Number of mics
    input clk_50mhz, // 50 MHz clock input
    input wire reset_n, // Input active-low reset button
    input wire in_valid_flip_n, // Input active-low in_valid toggle button
    input wire [mic_n-1:0] pdm_mic_input, // Stereo mic input arrays
    output wire pdm_mic_clk, // Clock to drive the microphones
    output wire [4:0] dout, // Output generated by the multiplexer
    output wire dout_clk, // Clock for dout
    // The following outputs are for debugging leds.
    output wire in_valid_n
);

// Debounce the input signals from buttons.
wire reset_n_db;
wire in_valid_flip_n_db;
button_debouncer_sim db_sim0(
    .clk(clk_50mhz),
    .pb_in(reset_n),
    .pb_out(reset_n_db)
);
button_debouncer_sim db_sim1(
    .clk(clk_50mhz),
    .pb_in(in_valid_flip_n),
    .pb_out(in_valid_flip_n_db)
);

// Generate lower frequency clocks using PLL.
wire clk_20mhz;
wire clk_2mhz;
wire clk_400khz;
pll_clock_generator pll_clock_generator0(
    .clk_clk(clk_50mhz),
    .reset_reset_n(reset_n_db),
    .clk_20mhz_clk(clk_20mhz),
    .clk_2mhz_clk(clk_2mhz),
    .clk_400khz_clk(clk_400khz)
);

// Logic for in_valid.
reg in_valid;
initial in_valid = 0;
reg [1:0] in_valid_flip_hist;
always @(posedge clk_2mhz) begin
    in_valid_flip_hist[1] <= in_valid_flip_hist[0];
    in_valid_flip_hist[0] <= ~in_valid_flip_n_db;
    if (~in_valid_flip_hist[1] && in_valid_flip_hist[0]) begin
        in_valid <= ~in_valid;
    end
    else begin
        in_valid <= in_valid;
    end
end

// Convert the pdm inputs from 1-bit to 2-bit. The inputs are synchronous so
// no synchronizers are needed.
reg [1:0] pdm_mic_input_2bit[mic_n-1:0];
integer i;
always @(posedge clk_2mhz) begin
    for (i = 0; i < mic_n; i = i+1) begin
        if (pdm_mic_input[i] == 1'b0) begin
            pdm_mic_input_2bit[i] <= 2'b11; // -1
        end
        else begin
            pdm_mic_input_2bit[i] <= 2'b01; // +1
        end
    end
end

wire filter_in_ready[mic_n-1:0];
wire [15:0] filter_out_data[mic_n-1:0];
wire filter_out_valid[mic_n-1:0];
wire [1:0] filter_out_error[mic_n-1:0];

combined_filter filter_inst[mic_n-1:0](
    .clk_clk(clk_2mhz),
    .reset_reset_n(reset_n_db),
    .av_st_in_error(2'b00),
    .av_st_in_valid(in_valid),
    .av_st_in_ready(filter_in_ready),
    .av_st_in_data(pdm_mic_input_2bit),
    .av_st_out_data(filter_out_data),
    .av_st_out_valid(filter_out_valid),
    .av_st_out_error(filter_out_error)
);

multiplexer mux_inst(
    .clk(clk_400khz),
    .in_data(filter_out_data),
    .out_data(dout)
);

assign pdm_mic_clk = clk_2mhz;
assign dout_clk = clk_400khz;
assign in_valid_n = ~in_valid;

endmodule


`timescale 1 us / 1 ns
module mic_array_top_sim_tb();

localparam mic_n = 2;

reg clk;
reg reset_n;
reg in_valid_flip_n;
reg [mic_n-1:0] pdm_mic_input;
wire pdm_mic_clk;
wire [4:0] dout;
wire dout_clk;
wire in_valid_n;

mic_array_top_sim #(mic_n) mic_array_top_sim_inst(
    .clk_50mhz(clk),
    .reset_n(reset_n),
    .in_valid_flip_n(in_valid_flip_n),
    .pdm_mic_input(pdm_mic_input),
    .pdm_mic_clk(pdm_mic_clk),
    .dout(dout),
    .dout_clk(dout_clk),
    .in_valid_n(in_valid_n)
);

// Set up the mics.
integer i;
initial begin
    for (i = 0; i < mic_n; i = i+1) begin
        pdm_mic_input[i] = 0;
    end
end
always @(posedge pdm_mic_clk) begin
    for (i = 0; i < mic_n; i = i+1) begin
        pdm_mic_input[i] = ~pdm_mic_input[i];
    end
end

// Set up clk.
localparam period = 0.02; // 0.02 us --- 50 MHz
initial clk = 0;
always #(period/2) clk = ~clk;

// Set up the rest signals.
initial begin
    reset_n = 1;
    in_valid_flip_n = 1;
    #2;
    reset_n = 0;
    #10;
    reset_n = 1;
    #10;
    in_valid_flip_n = 0;
    #10;
    in_valid_flip_n = 1;
    #1200;
    $stop;
end

endmodule

