// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vWjlj0mzNk+rqywp635eahC1NFzJayXDYzF4KQk8RnuhTdHzD+FGlXLBUqiZ2cxaCfqFBim5ip7K
5hgZIB3zCg5kZoRVsmNzpYJsrgddRcvx79fh+TwDXleoXv2MjtfCGGSX8+O5REGHOLGJGfBVBTw5
SjDFFx/sqGd6jduBrU9s4bK32rP1jkaSEkV5Z2ybHsRpfF15DKhV3zQx6uA9561rAZghA7K3D7z2
c5TGOynj3w/cjz26WyirWA+Qd8hTHQI0XIPWGHExh/kqsERKrY/ySnG8NUlPq+tbyAklQo9XHRNp
h/npzhio2QmHoM18fChTtX59iyhOv8Wl3kwtNg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 1984)
xFWVpmxmz95t2/3nKijHb7EgjInqfPrj6bQFhY+/rKgIouY3mKQUj48lt9TYPlAI1/I319edYszp
8/onfkY8r5Za5zp2ffFkeZKf6twnpVDchsBWbZH1Z7iwm6XH3misI70eeqw7D/UQ53guJ6VjeVV8
21fksESsI9K2vQhjBkJ1cuLevfWla9fZY4eq2vJUzFMfhqDrU4GP+x32Bb58067Ov7ISR6GVOGaJ
OaA4v0HXwfRDQ0zQ1DriuvFs9/AaRFI0Eb5FXDTuYyhReKj1BsFmxjB61DHmBWHtoEGRa4k0PkSd
cJEoa12KynNxaU7bBji8cG0Xqm86fAvfpxnzOUmVQaHzEXkIlU7KAxVO1YOhuwCez3s9Q1bGEpIm
Ibo9oG4FPM3coh4qvOX1Kb9EuYTvo8bSxgOyinVpqvMXIM0cDzAMPNrDWF60QSEjBnAzA21wbJNR
KsIez41IQegjA2JvudvzrwOggEVwLl5uS4Zosb33QitHrRFRo7dqL4O1/nROn7r6wfWQxTNqoB50
EiO2VxFG6q5KGaBwr0F/+Xe66ocF8JIq54vK/jmedfKHiPGjGK3tmGVE2EEmkq/y2ZpxHE4f4/Le
d3zapsTX6w2ru8uYxtu9xacF4rtJ3pMcRlJvxkMi1VFAugxBjAsY0ng87ko/DKljdIGFfk3zIN51
cTrZuVfsRKuSU4zocP6MmBarH+05gGbd6MkXS97QXjgfZN1wZe0nXY8pRQDhZ/NzCCj+Sag+fVTm
Mjp6JuM76AiecJiBbAIDWTpYYXMqMH0HQIXcwFrXbnQHJcceKwZzulOkgjIoArb0+7ByD0fCDTVe
4WDeHzy+pHvHcnMEwLu6rMJPP0hD/eVDxEtZcZAiXc7AJjy2Ku0PLzKFwe4enlFr7TUssWZMLfW2
N9mfFWZ5c4JH/r7ZTsi/U9rspGzkTsiWRORLT7fyvglJ+U2nkcG5LXn/iaEl4Pq+dclNVd4C9EzI
uxFxwTbtzCmrETMaZm4hGHCZJZ+bBzuMiSlpWvSBoMJNeD2erQs9+X9IyZEZpabrLJU/Nb9n2gxG
DdoDMi/A/CRy24xFgWcS4ozyzZ9p2HgGZHAFLb1NlB41s18JOoweQTCMw/FFyC2DL1i3TI3MBHce
wuCodhNijuBLBgVmmTODSRSRsKWHlYeahtnhPpq9+l2NQfdtv7fxG+vTc2Wm9ouZ+T2bDpokAuF+
ve4T7UgezeRSVf2TUOxHxmsrc3IcI/7MXfIG1ANL2h71M9y5bE5NlwjU7BUdFnv/Hm7wIQdFCitJ
ZEKCa+5K+sqPZIKV5PmdW/I+U4hwe4afmW5AklA2jZNU92HItDCByoTK4KTMBK++rgFWDEZWqPPw
SK5bklEd3nl/yobhHyi9bcvcIkA3xB9e8DIs3qCPplb0kVVLghC2uowwiJtRdtfCGmYszIkdTHT5
L6zYterVhNWjyi63z+2RCKwwWthEplWVEY4MhZfkSOHr6ho7SJtX/LfNmWy4rr42YUIG8Ir9BnE1
kEytmOuC5gq3SaPWJbo3/i5nAJiZ2/hZAS0o7f87Q/XSoxdX5op6+JXBMEOjmA/+sqfA/NMPQyLG
OlPoMqu0sz4Bjq5uhZqOlaQ26rxTVuvo1kjYZwq0Mxp0THPjBIOHBVPVkuy3YO70O/Z2uGVKqfM2
vmwlrrwsSEO+tHZNFGrtTQciEEDVBRGnoHdf4G/2Tm2t+Wxf1ohgqhBf1o+Ws24PxTlpxQr9lJIt
yatio9Spn6mpg/WAMzPP0AyLjhpd7g2jaxKcLikjB1tyStm59PrwrH8q9kxC2TpO7+xLW0+hEKLV
WQievfT9fB7XhqMakIOgQxGS2Z/OEvFCcCyak0KDHcsfv1tMxXM8f1LBy3MyN5vtJ66fbQIn6jKE
a/Nc1xijoR263OQr7QBFMIDNvwWVS0KwkY23YtgIAGLH9yHk2oR7xajo/ttpzh9GeqMKJ4s38jy+
9Is9/8uo1CxCMFlate/FuhTZBszYMCeuxG1mKyqGI/+M/u0lZXaicQPQBGo57v0OVBMHAOq2HPFM
W+HQeUPdaCaHrm5Nuz/uEug4MPYd2oo5rpVApcwqmT0f0gf+LQKD4Z5EqAyBMZehizhvu3aLBDyd
WiJ8+yzjBCx60Knq/TO+5rgQMAcm3Y1nboEhJ72T+lnoNWlBPV++y6rLT3KMoqnqqqiv2P8vlnT5
XDL18wz5fJuNiRULdDF1xHtkffB6nVs2CmykaowQ0Je5gEjdfpibs/5qDOnnll9UOyDScIJg9WM2
EgV9H3CRStfpEfRt3lBF7Kl3EYK+qFyZe1eILTp9S7ZJNPT25CzIbfb7cG1DxuLAaoU5d/UVGFzE
Y3uHS8NTw0bjhA+c6ziaK6XHdzzSdxf+5XNUA69Pp9hVSQCZEyIGjjHtLG7XL28F4yDlW3lhipM+
YKIOhpwpcR7T8FqXOVeXryvdsD9le03VXcu5Xe7TmCy7EpSIwIRH9ZXqTAAVBe01t0PTjihLKftH
GSuolfasj9Ln5dEZ/8oL4poDmY/4TqbAvzv97Fplt185MfKDu8vyj0iSfelkaFmMqlmJ06tQbt1k
YnznwpAnjKg4Flw7OckDTiu+TN26TrXdeG+JwO5XzqLzNiSTLGhIF8oK3ysMkw==
`pragma protect end_protected
