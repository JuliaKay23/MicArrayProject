
module oscillator (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
