// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:15 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QpOM7bN5fdcVJnqvbDxcfZN9+sjFpfA/vXuBiTsRAqscQYePuO99n2gym4llbV7r
E3IalqFPcabisAYAJphSsLupBmNcg1K7tPmMJtjsp6ryu3DyGBnXEOSHEaCKBwn8
4GErG7pu4aFSBnpKkNSS3YhwAVBc6UKh4XLnozet7A4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21296)
Jq//FNfrtPiO711Y/GLCriMNLjUD1elxJs/0UaRYcRc+Y0ynbK8DYTbkjSbrFcqw
Z1NwIpveFCH29S4glWM2LqqP0v4m5R7ROdQVpQSHI9yopCk9+6sO4gZ+aMppJ1NJ
oJgXoh6Z/qtOFdcjq7f9uceAsWvN/lzgL5HFt8hj6HzAUELbxsV58JakpPl5+KsO
U0rahXrgrciv7K/bMdFVdiSvvIf5F8e2lbEXFNFqOUL9AjzznyLTw6fWF6C6nyb8
kwVqz2jfp64L9QP2qOcYAqYtawv0Ifoa55YVLKNvH5aVNSn6bDCWkauBAjDcJK85
1YtprXyyqBNUQ26/a6dJGRJrAm0V0jny3nSNrAi6I/ICu1Ai+ATtjd5StiOjZhYu
wBnzCMA7embPsHVy4Jk4JspTyxyIX9DwidLCwSd3QOaXzMlxWzM4Nj/HVGcwXATQ
5M6eP6YqqpgC2llKo+gemju5a8rZlWfIgazFs3Pf5b013QDrd1ST+JWocvGsOy5Z
4NxY9A5DijYtS+YsuTZNlGAcE2aWlpnHsNOswGaNYn3ntP2Z23F/fyuFOkE9EdC/
9Ydd+1hrd0Ke+KUYW7XNRWoX5lIbqKZkkf5H8yTqruiHMi04QWxKGxhsOwdIYnaU
SWvnJz+p5E5W5/yuSUeAhAZHJk04R1QpdVoHJ1GYg/PVPcUH3mZy4x53/44l4lPA
ykCpbnNwGpBu+4VJdtKaVMAJnwdRfD+Ott2eP3eYNZl/E7TmxfYBZ3gESCoO2EEN
UzXHdLyxSLm9oDKgOlS5Yidas5+9qA0eHuYk3N1hrZMkk930YP/809+1e2X7vX0J
2Y3RUNlpGn7ZcFdNFFkoMDF7k+Q1h4+04nEpBNJBi/f1rJDvfGqdQuP8rLPZnKHe
HQq8QHLvEtonli4kq2/zdAKejQ9lIBqudJ2xO8dSjJS/uradQSdEBFp5EWdshk1Q
nXSh77CFDOhjTzZLe/rU3FQp5XxQReFh30UHvDhBj9zFVol3sL6giqzYPGAlBork
AnqrwU3QpqaSEZpQtcK7xsSGQNu4xIkackkC7r9PBqU0FL/izPh3sc3NDLesQcZs
3ChbOzsUvk1yQ5k1UBe3lS0OIjiAQLM1wSyKmrkGf2YS7RWmXx3QGUUbxeMvOZKS
0jfGzBHC1++/qzivIUkT8s2uB6H6e9n+159TbaFlq/5WXu8+I971qbIVmN76Zs2a
39tsfvFC/wmUGVrMp2GjicO6nrj9JHCyeHHSBLSzq7dtMD6wj0+G9ysaLHQIqYYe
6OVLJtv3ohsQuU4JgzbHC4nYUQK8F9jrKBsNQQSDTFCtaTnOG25rNFYXXIkW0Z4C
x1GTxKhGkNLDOF2xpE3KaB6+0fVvpS4ulDU3KvzhL6r6lCvLcmQVZd286X0nG6OG
twDlJruCxx9c4Tj4KSpd0q6zbWDcirVGl8ks8JgGbaiYhmIIfeO0PW9J9QCIU4oA
/BOQoEqJiFsA5y0RzcOzF7GoXwv2hp9j4hiRcai2y7RD7Q5QTMecJzeda6gWQ/iz
cht5G8q+GJiXnNDz2Ex2mm1RbGLABuF6ZNJpHPomSU+ybuD7awHnzsMsBl9f5+Py
Yg43aR0IglY7q6uOaL9EFKyvtSzGZXLhJLLW764UFcE4QbXqiAjn1n+A/rvIN/Jx
6cph4ptJs2o+aOIO4AZ4q9lNTM5rtm6lHVmOa06Lf7QyEasKgP0jNf8k8y3Pse7s
YAnzLPvzSlDCwmKYG5R7M/wNwxPSUgGyiHIkyrNoZvse1KPElh5DcT9DEv+UiJ3T
hjnSez4yfDb7CUjN3LCSp1zAYujqRBGi51QSP+Ke6zzlEts7Gi5RrzTlUWBg1w1B
vTY0rJ75lzhd/z+vZrSmsD+KK8rW8kMcP4w3FlnVxF0Ij+tJ2HrcoB8+2t1scFKa
mN3zLVp7772hDQiq2IpoKX3P6KqfAK6b5ZOP4CBXdRVNPyj3c/RsfJQ6LPIqG2bz
oeVxZapyW7pqtUi1Ob5HF8V4dhZgdV19KDDVwiWKcd1IKKhpLgrtyXrRVqlsg87W
zPGqsQzQczS0uob5uIzwlgyOpi2ckM/ZgqHmMGNBELv/6TuTmKJZlr3tcfWUeAVs
gLPPO1syXcCrzj+Oqyg76llzhAGhWEIa2gP57YpQ15sTbUu7YYZRs8gXYmyU5VFn
447pzn81BuN2cX8ZfqBACxFthqXjAvebbHwQrS2xYLo4OFmtcZTPervMvdzYa0Nz
zcEWo2mxAZqETh4ijqAMYO8PE1W8vkz0MHhhs8Ovf0RULn+v/WdSRhyK4rRZiWCJ
ulMnDVV8eC0SO1TqnUkH+lAi67dHXxtsu5C+tcggJByqyTgrAYWjvbUYoFKyHixT
94+gaTNxTRrVWMOm368dQljc4aamyuSt4iMhRneA/C/ikVofaYE+qrtujVUQYF4P
MQdOyh3BRVI2gnnGbqfcrxHSu4sHg2d4KK72Cj1shL8PFBMhXloxqu3XUru+sJeE
6HE8KLP6661rHm7HZYzXetCRvonr35iS/biaOXcFJ89yKiTlzMxKzzl2DahfGYvF
t2nFq9A7TIMepX1YZ3HbpmHs5MI0TJ6cY3FPhCP4RaRPkXO0p+nHmUecWlOk1UH+
E50D3sZsQ7gdlWqWobjl7HuS365HJ7A+O1kHC/kTPbtu+BdUgn7DrW8Uz19tTUC3
CHwUOQ77Mrq0h91p1YK4WaWdFfwBEPlVc8keBs/pxbBzicY4Ggur3TLuhXDI317X
kOnKoIrXXGys+HNXou1eBOQBW145iqmbomqCWbDZBLOwvQG8UIM964fynvQbhYgD
1lyQzvFe92j+9Ii5onyHrbBD/D21cAcPT7Ns0Q1kpcfOHBcVrl3p+z2MuH5vgEKv
eM2FvEDrAX8w6r5a7q6jE7jeRVmGgnIecZdkuN5VUICzDUKwrox8bDWjIkFbcsAF
t63eiCHBTQjOHkyvy+Ivwk61CcaTGm93ZMGiN7Xj91Bh2jYX2yWpUFMJ+4t9yHQN
bXzchosp/eBiD8cP3P6Y5DHVWwTElGgx3NMCAgOF9UUb9Q0hNT29s61ZrFjSEc9k
qVfOJjjH2/83AzN2bjBWtSP5Wi6toB76TuJs6BH6pwPo9yu2A7fHttkhE4tLFmy+
QnZ06LDjZ8AJecRIkz3eSXGjWckcIdXALRJqGDEYTjD37+JZW+klpGbuBNWHcrQc
ZSFJWlLVuwWoSTND2RQu+DWH5evWePqRY7kIGmQ9cafRQh/Pd5BW8YDBO/Agm31T
Xgg6eHMSmKR/iqpeBdmaGjmXNfb00DPuNRQm3XlXLHDu5jUMfBLPKxMcAZWIDxYg
VIJNstJPbG4wpHYbpe3J35BTrRLGUkwZC8tbXA9++qDQNQMxo4vApjc45UtakkQH
/nrcVQiAIJM+w+Fxoy1N+3EpVaiIeSrMuFiZ73ApVXiBqheNxZDPfXgTsHV9/6gT
RX2FPwaEKMFO+NeRlxAJ+5LTKKLpNWz3kaUgy8k0Cjgf34W1PxC8pbixfvABJOfL
9Z5jNVOUUut68rDC4p5RvphV4hMS05BUpoWcGmL0bJuxhUllBZBQYB21VBJ03nQ+
MswxKpS/Y0Eifud0OX+gflcvCCzoGPrveJZgpOkqPJxWX8JG4OLofR7nJv6hH8Ok
zEaPrbngbF0n+2aRtZFjKWm9HhbY5lNPpFaXseNrxXiu+h3+PSj6IRMaVrX3Kvd6
TrCgFLhFVl3np+/P5rgy4iP+r+UL2aeT+HuaStnksTlDuN5bfyIgyPPa1cQvQGB3
NHDY4pQ6Ghxsb9jSi2QSCXjbvroYnRfvvwyjoMFJV8QtFnAynfhTf2aFYhw02Xap
fO8ZstiFB4z2KSzZOZBdypOKNFOSjE4BINyKIPzYxHBPJDRewN5qGk3d1HVCwqdM
2KIJPBKTohGHFTltqt/7Abpd6q1gaVLtPoPtZhZuzs4gxOJCZrNsKApn30c2T1K1
R32DYBWzA7uDb8ZYxKMg27Qgc5mFesW8vDkFp3x6Lm0bbnPWWjiCjr1L7Ic5O8EU
SuEYKOvAXqegQTukXWvtBRc6oKJuW8Cjwd7+hwBpsf6AG9maWsdSYbIUkqVyv/Re
BK+dv+C1CySxgcp2l+bA0y6rOxif482FMJHFOlHVuBPWvjDxOv8gfkQOHDwRzfa/
5nuzxuHUv1LpmEpzCyw89HsWE/E99xulVCLt1S+C3u0bSzXpxjo14cWfpUsH/ufD
H4tYssko+C/2KOzr/Xf1c5vs3WjWK6b0APG/KOo7dITB+yTpZRRoKrARnEw978cD
uDoZsvtzZNIWvMtVuxkxrKlbcCbVRzd2HZWF67HAs4XPtXvfTv/zZJZYeVxNeVcq
RJmHMsRObGy/ARFJMCEcTlnImdv4YdMi5gMrvTzJesolkV6jrUooq86xuNizSWFk
Rd1M9f3cqubWbAcVir8KCKdnhSEbp2qMIMgac+8BgDAaEcKDMn3Snz8WmqDqC1Io
RSrG/8KNhBm5mxPpuBCe4S69LB2jUz/8LjfkyZnxPEgVM9r8BIRmoMrfC+m3bbQx
pPd23wvYecxK5jzgDparMSUuZk5957tkw+v1F6WYTnBFNWba38zytqXYy0ywHMHJ
m3oSRyFpvrecps4qgqlWDONsSwv+mPglLuMqNGxw6y/RRh+EUZfB/fKtgnBLUqTS
1AiyPmEgj99DKwpufeKZiwa8Hsi/vnTYWb9OxP/5ZikO02jmRBzbLnjp56GKwPGb
kAuoatmYgAPrGXEcqLT+YgBMz/elL1Gk0v0sOUcoctBH4NAfZ2uRB5UA9YQMxdU7
8MdH+YHtJR+FvfxdrVHDLNFOjyJtjeuRpE9/iTg9sgoyZ3r9Z0bQCuXodmD69GZg
ksNUD+V14wXH/zo/Y0hbj08e61zkNC8Lg7/VR6cbgU37eMHoCIBKU4XrZ8PHXTBs
BaCRObuSrQronq8rkeG74Mw+EFlGw7ssWraEFBVyW81/KZmxgOwF7h+rf6IVQ6Ou
zP5MPUnt2fKnnGEt9EVwSmK9CCRZeA7Foodw6qlYGVcBrzD2TG0k3AQz5ds1cCcy
dwcfJYz4msqcQs3WmygmKpB77tVrHuF42uKBMWi2Y8jJn1+Lg44a/Eb6tOdF2s96
IsAJLs4FGoAmLGuKcSM0l3sAGiPm6npPsfP1qP0em1OeSqb5p3QG1ROeGaDNUExN
tb0FoqXMuvbNRmPRNjZKR6hwiK3H79FEO8fapNY3bCZTYba73wIdQWuGrC/q9kY4
SOIDBDEt0HXuhNjex7MGQtWeRajF5+GreB6JQ7I//qgYslbNXLi9rxVsyOv87NYR
NB852NKaBb40ACzzAZs1WNh9AHbCF5uPsKWN+77MRKYP/bYvsG54Q5uG+elIIAWY
tmacLsihRvCWzQoS0n6snK9VqdQUZaNu45Ruk7XJVbUNAxn+GYqSawjkBqk/hYg0
VpXU829/EXBG9W0oGH7qV2Q0iz1KfCGq+k7OFO50FfYbSzE8bnhBMdMMgibGyLRv
3NwwDPCYNZWqCxRd8Y5eSiws9UCu20r9c8YqJagLPQD7MdARA1Iu5MWJuqW10TsV
hXfMgMzTzah8jU3UHGFfbGMBVp0vPnAc4+223twGQNMGuhO1VsYzD+FcAn1VyjCE
UetGDnLXbtYVdq1LaQKR5vqzSc77DDpwsph9PQg2FY9DdGg4xEzi7Ly4XC1a3zY5
BoBXga8fyF2M0viMVt4nWngvc5vboLuQJDeAfMqyMgt7psADJnJkfeb+6gv6zg1i
ss1PwkUB+vCdJy3U+/XbQ7ro7delpHr/kCYgYroKOAPI3JD/tFqNoXCDd+kNRUjj
l3buUoytz6PklaNMRwAy2MuyD1MCxeQbTWDa6dNVwZJ8vhtDsIovc0SLulwtn36H
HFAJEv0NQVkE64UMGh6BX2215y6wNzzry/LSKDOk9Bj4khNB1sTJ2u2XPVLZWhiQ
OC6PGREKeNHBLMI/8AO6UZjiOi/4VnDkxKLgUuoY0nNa7n7NS3c/tFr4Kxhc2/et
MXZblt3+KY+xxggG9GkEEYBUnTKhCCW8NrMTMCyyBlTR85d09gSmmumacv4lteOA
Ky1jhn0SIEOQ+90SHvOT7y6kBbWq3iK3QMDOP4tSSdnxURkrQuAohw832Z2o0QTf
+WDJX5IVlW5A1Nn0tt2KOYzGFnf8jXFJW+Xwuq5i3Am1m5ST2vzAC1ig9stggQMD
NfbFFzdppZLq3t4Gi/AWSXeFMQJgMWlhR35zxwxFz3R7e7ZjYIrMO58gjn8teN+W
2YaqqY/Rofj7ZeqTfR1qAjiGuSMt0lYi4am3FsxDy7B/h+7HZ6qH9vlgPQTBJUGO
BdFvZhi26VVMYwFh35c2NSFRvhbTdgkKPlECEI4OWwOVmAl0cuWhpegAYfvBVEMb
wQJsjWaRjUYOqXlCEnekM1dBKi0WzCcxj2mpz3Q5I9acnB/LI5H361NiFpVySuE/
DDAj4CeKA4/qmPFVQxqNZL2sACXrBSHK9MnFidh7I6DBdTXKcLOJuxm+eIol6iJB
0D10bsTlT0ApAxXjdOWLDzsJvdcMr87QA+N6ak72hQKwBiW3JdDtV4bYKkjM4Ana
BHun6/8qIgnA0bY0CCdkQuJl2Bx05l5fR4rFf9WDAoHNHSjS1qQSUU2f1WAXBUF0
VGnbYP/lHxmcJai/kbSwzEyE3Aq1dKrT67amG3yjS/g3ok1EKgFBUQ10gU7F8+NU
bEFw4fZBaAVwQfBqF7moNp9kKrvk3Viv62ViCILD/jZBCQpEMRobbn1/CsWYl5FB
vp7YwWGdJEAJeqHpKb3hWRA5igjJF9PCuAWjOq35Dq2/LCjPW71C/RK9yG9BxREM
XFX2t6FNHQEuru6TDXsmhhLRV+zqTFUKwE6oxNzUXkVPCLpAOOeNPGnsXHBQODAK
0tzT6s5mJSXzd0fRWbGydayY0jp+kzjPufVgdeDdU15p3kj5t3Kgv7gD6YgHJ5KA
SOC6kDAI/Bn+cWU0ovAdF8j6+BxyA81yKc85UV98AzKZKkBvTOl7qwvAUP4l4jYu
e8SP9gp9bxr2fnoKSbMmd6KyNKuDT7cgBym/vlJah23TNBMl56Zh638cfp8Ishrm
uFVm7bZl80XCpM54auR++KI34ZrRcvl9NQ3AfldsJNZ1Uo0kSeeSd437AWjfs/VK
L/Zt5y4DPB7s2IjNcj0WoeKU+p8eNz8fN9B+2VxHZ8CyjczUXOlFu75oQ2ulTvZ7
LYQd/exXaAuIwc0DuQheiqpXuv56WfE1qGXb6iuLNnDKa6S9dDQSdUSgiL1jOYgn
yKcqDz5vLCTjUfPLBJ5GooGJ/NflQn/7Vfy+e5oCv+yyGjGjAw2XcM/hZ0EKYGJv
pSCYX7Ny/LUdwboy7S+NgZDPTaDVShuieetFdtfSHeNOiI+z+wk78dI85LhWT9nG
HKNhClTbrbvNqZw4C2mqZe2VdHr/LpNenqgSmUyT/jG9B9gjvNXc0g8pddtPDLN0
fBW33leXkNQQDtww9I+xibiPpP/nJaP9wfy6jDQ99H5ojgEC3bisl9jPMenqWh7F
cHbkUfqzJZTyysG/UUjqj4hskN4LIv/I37W36GSrJ1ek86v4JckI7n9/KBxsQwwS
tfgAoyqtpDzCpfEepYPX+1FFOVEDSmWCgsLvZmU3C2XBR69Ctx4sAFjTES9aiehR
5t0kraLBF3j0cwCNVYncOfdIyast2FFQdQ/1KQsSFtbbq4tUbA147fHDc3keFr7c
E4A5+wgyCSG1/QDBGLFxEjP+j7VkUXPK+0agdZ5omveFFovBjGqOUlNrfilXb3LX
+BCVpAn76epZXc4nE0mGXjQY0ZVLIENjy4mINimp63l7PnnOPVOuwhMv9hdOlnrb
Vc8BuUPCZxeZwDwAxBQUzIIuJ/34kE+QA6fBZ06TpySJ4GtCOgapc8lIVldBFYm2
nF1tgWOoNa/ZvpL6uotNijFyKudea946qIWDeOODPlU0DPxtWHCk5e5Rkv7r/0Es
QynDKOdJAhUUHuVsY63qgCPmOfTPoPGlgUt5gQmt3leGQ4wysSeG/lNT1PtK93fS
NCP6pcK7+vau3U2VA/Ype1P/oMPykAkObSwH3elxyeiDIG5ehV2stmCu59q7fe5k
nEpXKVqUV5lSA8IKbMFsYykUn9gwKDtaVQEq1u9oHwMMeR8cmJZEW5pzynlQ8ONe
ZrQGE/nKX3sH8iQrtuARHVl3ylTcJPR42SqggeCwUEDpJcs6IfOwIKmLhA+nvbNN
940CfDi3996SryV+9x1Zxw05D8kARmuYhy+CCvq4KDT7T6mR+2bSPDAOdAAuvPG6
WXiCjLX17gQKq9YvAdGZcNrIWnlN48uu0MQKJZbl5p7lb6Cyt2dgipSFLfqs4QF1
jii+9Jj9KtHmKcDtShPWXQ8I2U3n17ShZEeMefcfOfjwYlX9pDa1r1vzXI12tysv
1f7fn41BlFouREx02U9F2h3vIC11ddbGrLj7PYanHhFN868Q0SEC/KNSHziOfZXb
RznAjaeuOpds4ncxnErPUNmLaG8KJY/NSnpKaLaK9/znBhXyvlpfkpBnFreC5BMf
4WfPAOEqqqBmjj7UL7og2r66UAbYZKff0C1y6VTs0q8luEopzpEJLSJDNetloonV
4cIpp+dGK5K77VLMz5/JJgMfSPkBaeUv3xA0ivzk/AvXtWqcQeMgm+mdVjwk+uJ/
limbQZsPFRaCDbC422yY0Z/bZGn6siiVcduc4fsPsKt3T4xhzJXcYF1RuT2KPgrW
EY5NoymqV27WDgdcq3OnZ3gx6+WOFB43V5cRQ2kxyF5IKHrU2f/1ENDZ7TZHzwjL
HyhBncLVD8PfQLSOPQyF/+BP797IsYRhL0omT/qvFEqq8gdnEtOKsO1+ibWuLwHK
O4XPVXU2eVkvHvdr93X+4MCfW5l26B8M9UJN05jX9bfwUzplAYrxNMib5dWsP7+T
2GwIpWR4NNV0jJQJCMO0O665oxNB1DYgNAXIqgqFFT3DtRpH0Qld4UUliSSRXO63
syjX9lhRHdf83bRS/3TdeTu/VfCSa/pn1ctCsG/dMc0O4OR0BHTrqeaNXnPlf3g5
pNbqLjigV5bJcHOhLKLbz1juB1xP87uOABGMAX20ylHXP6vYzR+tLCMPQ3aY37UX
IboYnqQa/G+sfKIb5dBswZ+HBhR9peHXVbioOpZVr4wBr4J2vdQIQFWR/nShlLKW
BzlENDgrR6DJZAlMK1Bkbyh3ue1rmEDVJ1w6Kml6sdIYEcVHIBcDSQZeYdTc+glL
zAvYmU6DSvXSDeY9vTssG3Yx8nDyCqTfig0cjJei+9BH4rqUsOYoIAFBEMF/KisV
+qbbhQlD2gjsvOctklnz50KVXNnVrGUfar5dLvvHVo+fSbjlGGdFWkAhciW1AUUb
Ytu007YPJhWDmeByyXzdh9Mn3aSRL8A4EnjQoyrnLzD+aMs7b/Gpisaj2/MUf+5e
xqhd3jBfcqRi3s1n62nZ7V6GhV46C7f9o7mc7DOPIc6zenvWlTwUpACYd64ESVxu
Wzq8PircQM49cEKwpx2yqaDYFUosr+C8mxwy/l22ALsQ97ZW0vMrbHlKnwZt/8Ac
jONV3Ar2NWPQZsXb63BT6lV63/sh3Yqoj7zFuCqYlg+iCdTgw67a9RvUzBIgaFJ6
MdaZCz84Iv/79bAhVNJk8cWtRSXZOEESHcigPJRL5CihgCNnxoGS0a9wlvX+e+2E
1jj4lERESI7FMusf5It/ohh6vyhXuu2J7WvBvUlgpaYo4VXH+SNn8ykvz6pggasr
P9xeTDob6VCffhJ927oNCnhd1LFjleUEm3PRCTjJnqjyfRBcXTlhArMbNDoKnw8N
6DEWWcZPRi89BJ/IdjhTfWEKfWLtGZgXdpdzWJrgm/Sw/W29tyD53XX8EYwqPr2w
1V0WAyNNIvKPz5vMin7rxU+Mim+Zzm8ck1WlZBCdVGSaLMRHFi3UWdb04gJtDUWZ
ntgcnkA5MaezWIMjh6P3+7U+TWsKejbrGJa/FyRWNYo0s5OxGAGivyY4ws2F86d+
gzOiLZr3KJOa3bm1JBdWq7P5x4Sl7B9QBz0MLa2PMQQcxZuzZDiI7ornKyTn0WjD
JtPkvA1YGjW7lFHdE+AofnrSSy4A28zyr6yba0+RPy2aEzqFVDwk6N5tCjkaZOrd
NcYBWPgYWQeCAbcLN2kloL1zTJheX/81iwfSbm6XNqosk/XYx8HTKDgeL2jfhwew
bGt+B/bZV5kza2YJSl+veXZME/UQraBA+ItZYdE9oEM3Vc3ajqX1gmgVEK9CXwH7
k/B5muwMon0RGgZQStPBhmFVyBvY1grfTCHEC6+t99QV2JFbFy6IZLozYHQdSpts
Uttuapk3aYeu0G/mNzA88JSBmLbaQB145c9cRsexx4SrVeQsw/hEPhrQZXMjBt44
0w90NGIZ9GMpZVwT/W4uFm0wC9HXAVGDKf0xS2U4BpcQrXjca3s/dhsAv5FWeEUE
K/D9usGljA8T5pbU8tQis6owjt6Hjr4Y+uw2zToUkBOtcF7NRYiE19WJtiEz+qs1
+aHaj1ngMtdtb2AHInKLRFojDyrP26wLoUdIiN1TKFsV6IAYiFG5ZXgu1kTSVlEp
D+XBsn1nx65HYPg4MsKlCcaZ2hHZqjBRl3CnO37dAUf++X8qO+y/jWXP6etBtezd
Pkgf7plUCR1ksOmsz/Yjz3fbIfeng7k/UWJQF/QNG55m2/efWpj1n9QvDc3Q0zKe
hS9Nh4De0iZ9cIixtZBL3x3fjlxDaxGo7maIDtbTZyO5rK403n/RpiwiBK2AWV1I
OvfS1Ynz1m8H9x2O4Yo23r/GCxJ4fKyIdWdtBgKM1BBCFbLXDvpQIsb5BEFBZhD+
3H506psfeM5L7evlLicYWj5fhzdFfPuiWDLr30owEr1h+O1lW08PqsnAZPkVeWX+
9ENGeeqHIq3U5cscozLOHRC2ykcDLQIh/zKCZtp/YjL+0THp1YT8TVM9t7tkaL5e
ofCp3t5Igam+wQtPf3BLJpAlqHfDZjt4jJHDCIBIj3utnB4ONYYA+iO7l86JLNno
tz6mEwwWnH0qgTt1wCXu+hsGiIgHHhnMC7T5vlw8m2aubZp5FHWTBHQ9N6Y9r0yr
Ne0GwL9YLgDs4/YCLYJVDFWPq7ExzhontAWee82DR4aNx6RU01xcsF79VvO6SG7W
4/Pptx1qhZTpZFI2xK9jleKYOx32bRm0vjz/0HsUabJVFDmxMmbDKJHXkZzA9u+i
LH/LGmEjKQYU93brnX2nVVnTaIVxcZTf4Wv/LP8Dwq7NAFU+LuMYnDirFXEbQ5Bs
VrZa+MyAx4KSY1q3kKwKFYlvQ/6FgmdZSB8i+tYQ7ASq1wqitmSpe+ls3kzpUrM4
dpsC9w0JD55GzajhAhnjM5yrfcudZpMYMI7DkusAI2YCgpqHXoI0jlqd1sfiOqj/
VBCnOMGsQYjpIBirnSZLxGp4lYJ0Oowq/v6t4Iq9smAieT9DYjf4ZvB5MsEHyRLA
Fpbjc93UjeUVOd9kyljFbrVSILzxXSIsNnXhMy5v2QPl5/ZITEetEU/qcr6uumRX
KxopNs1ll1wQzFv2w8JD+ISJuU1h8r3GPBsrssD7xJv9I2P+2t7zGe5U03bKn0Lu
z0dZlDZ2TK+UrTKQ6OJGhTdHWNqmTlzdDZa3YO2H9t01+MIfWk+F0qHyicLxqh/P
xuDwOvi5hrinWBMckmWEl+7XHdz4HPbQn68yy+qlmBIOVA3vItxS2dBR+RR9PeFt
dkWSJOXC01rNjKOoxcqn14g6smQMFdzcMLlddKyUqibjZPyyWYpUqlJc9RvK+s8F
3+elsp8HYERJ3QsGf/ywEqpBZWdjQSGZ7pBuGOeMuLZue8rvS9zwUYacICjgPeuu
axPFkj9ib7z5yRL350YMqg6ZsmdfcXJ7fVde9M8HN2+eaTeywL7s5PYelNiOrXz9
4yS0BdKO/1GIG3BktXD2MphfxCCdyWiGFZSH8Q69PWl5Dh4bErU8BcVHvvarktCT
JFqmmj/d4kCDxObpuOlPNyoBmKAkX+C2vWsuRIqj6Wgoc2L3YCKm4uC4rmWNNNrW
pwDZbXMYscRjleekpuPKzfxp7BO7p5fvYo96mIQ4+BUrFFFi8b0zCp9S55FWTHq3
CjvYIuOQ+0Q1OxwVe6l7qwibW/ItEL0kLGYAk8lf1wEPSHhrlOtvEX2OdFaabOFr
pjW9WoU9lK3VsSL1u9CqSM/ddwzBCVp7BbPP1eWVcVxCiFsbNjb+D7og5FMAuNhS
xChEdW2WyvIgPgJvqs6auGR86iQ8CbhKiQjIbZzWHzrIw8PxegfQFDJh3kWqFefT
Xx1Glk0HWUHgEum5Ic3nlTzswduraE58jNkIlJcM2KpF5psBoZQNSwGMAoQi7R5l
f82kAUEwU0/WtFOA/91D7TmYFMtotEPfQZbVjZvnwaOxIBISgX5sy0EXZG0pB01H
3a6qAHpt/Tw28yOXB31y9Y5DAaTAWmIKTo11C8mQ+I9UYXh4hMejetqW/0Vp0/Pc
347+QSnmCqDVJuBu2ui1iN94vXHckCAkQvjAtpkgZ4Zqv8NVsLcouzdBvDHMHGno
8PCHL4jwQ9h0E+ZDp9p7XzkBZecIyVdeZZ+VIrIuHZGEZpXik01P6RRUcT5t3CfG
qKm6wnB8W/7jFOGsK442xKGnh3vMt5/KOZkOSZraZDVIq7kwWeWBjOPVsbxQpLBg
ycOzOkXjsP+kxX5hmejZht2tW4Z3KpQVOaG31keK6e5IDjsmxtEAz9+G52qw6lZB
JoKDRsYQiQkZnQjGqZicg8VrwZ9ycJmGr1qmxBddcr7CJFS5xFV2luLSL/2HwKlg
RRHgqwhHyrXG6xi5P3VmrrjUQ/NXLrLpU/UVPrb/LbGsAA8SIM4BKrYmUcEj0+AL
q8TeecE2H1nLBjf4VlA7ylO1lm44nuXG7XGvMpc1HVgsnZ7+T8kJDFjccThyUGWh
vw4MSFzjdlo6Iiud0GFX7I3tz4DlDv9w7coiCb9sr918jbOhT0Q/IbjDERGsFACK
juQlCAwfvuT10DfG2Jp5jjBrFStWmMs56J/R98ZDQkrL8wII1lUGNybJKHq97mxP
gky0u1upmVxhELqQInPS1YmOjslRoYUzktbVTEds/53YmZwSlPYb3nOE2wbhZ33e
JbuCjATHdPHx8d5Vdr12OiK7WCIHBKCrlaRcFQN0udNyP9qtAYOLy2e7JLfT7q5B
TbE9xxYAVXC1mMbffgt6pBc4RmDHM1U+Rv85aPrx9roag7Gcx/ODqMRtnKrJ3XrM
Kx/sP1Xz2DlOrMUGaoQqDyFHARz/sGAjP4nVwEuJCjQeVh5JQzJZfBtLKYM08ZNF
cJEONy4RoW7+6rR/CGmfkhEnnrVDh/R8kt2DSuPMRbjV9s3p0SuvRFgA4EZq4ViQ
61X6gi0dR4dz7NEF3kO5EvPMiQgkXgjKNoL6PfSgOPWzLMEsEOj6IUnf8cXqPe1w
YZuaE3eAsAQzA3wfdENhILIHHeLshazoRM6eKzVkG5Pq3rcnd84ycvcpDxpdH8Se
LUG07Zc5zpKBjdyMDCY6GKKcKmaZ8PD3UxzQsG8TahPmEianLHBalpQAmVvZAX7d
ur1K0Ex8fmYZWiMo++uA5HrWotr3FiQC3xKDQRPMfKdhNjVSZlEClSHTOcm4feB6
AhhJxDFEpN0/pVvGfTNp8cLZFuyWa0nzevrmkbJZdQ4nbDxVOuQVFH66is+U3qU1
A7AGzUuBSI6OvERSglCyHOeAxyyXyKJsIIFPF02nIEw5mtbtdOF3hTmnZWKrF7eV
f1IwLYFSDUJgxJVZvcubhTxlBlce6aWCLh3xw8tqNCY+arnybURg6UgzyUMRQQc3
fZX4W9RU8n6A5sEs+q7s+JqYr4PTH+q0Osk6Ndi/6FIcdczPAMPzoh4fsvCZHrc8
3PiQT4nTsFzOa9R+y3br5fFq9CIbqVpNxNQE9tArNTOVtoyuik8kfWDlmjXKgoER
fPaTaKjmzYxohdw1bbSsJHdQ2C8ZilsPlA3giUCygJ8/7cBv6OuoBdxNT91ODZcb
Df8h4lA3v9KdBNYZGR5vST6mhOSv/j3Pu6+CcE8r8hlbWY2sBNb1ctaC0B1HgqYF
CWEeXI2ianL4QAXRqT+4hVzl2+iJMFQQ6o0ziP39M9vT6N3JlCDW4WyaSwyjqOnL
KTCyBokabrmB2A37p0WdUo2hPwlBQP7fgz5TOdGl9PgFumG/MhayqY3QSjcSu63h
XTnP8tBmCN+HwBP7A6UjajjkLW+7PdPp6yJb4I7NQxICrPk4E5ja3xeRmQmmQswU
vXl6zm+uBZ/kYurIF4cNHi9GmR6pO3aa6dTBIgX/Y+NFFgWoxPbqBamGuFeCmVUo
4TdtxUU1m9OV0JCZpGGxQVSNZLMXqby7cxzGJvkC065lAarN0NqK5n3hQ1thX39P
jf0kLuXfKOXyImNyTFTBDGyd4uueQ8OofMPBlkqzzINo1khxfRIox8OPpDeQVE3k
PKRjlP5nK2qZi9+UPxBS4Rf2EE9mDV01QdT2EmQ6M7uZTuTMY+aUpfd2197WJLIN
JUgSfU5EV2fybIPxLiggAGDwBXXi8eEo83IlUzCwI+m7aGjdZcoHtwuRLDDWPQL5
w6sgMYN2fvIbs8kB/Ql9Q2JEaRKJ2kmn0PEoyE1C6md315U2bc5oNj1u6ts9CNMI
T8gltGw0ffk9eRTT4MP0tEUXhwG4Dz9NOdv/5whdE8UpO5Sq4URnPKD3WFG0PSin
abSI/9agODYkbJ8+2N5JMbPoaCkdN8TPIxVqLNe4xrkzgmRIxS8hhG8ygAov18C4
aDwa+kDRCWkGB/OD1JlRVXtppJ1oAN5mn57tiMIYgQeRYK0i4z8OAYwC1k3BzNVq
Txqgy6tYbUaDk+Ev8hDL1cST3B0/lVOj8QQr4H65iYHap6NlsuYV5mGwW7Gh2Z7D
pGxgL/o/5JMzlaSosfOoqMebpPoW0YH9FoEvELCMQjchnyw2jQjXR4vuS7BsoYLy
7rs6m4RGQPA8TN9r3p5iMwAJnNRPE/wgbmRym1qKGU7j1S9/7Go6J54YkHhPk78g
WKWHu734ivhy60QPxUqHfdubJbrOmFaQtAJR8NU3Svr//stX655RJA+1t0bDru17
mjJd2kwpbwKGX/1powitYacdJHf+0mbCzLJ0zEIldVECMZyue9LN8of1Hj4/3GwE
Ymt96ArzGh5W+e4fwd0E+xtrry7PmdZi3pGArdGNMcOvreCHPLmyy460qyTXgAra
bp15aueDNwpPE54fDnIjCSCLnNWClQGIEBfnkWTB9zHkIJZkhOAhp1Ez9HkS79+h
uJ849sbW35G1KSBDb+Ry20f/nU4D/JzLhDkYQ68xMbp0f+nHeuYn2kWccL/vIi3+
eecq76n0DcRB93geJyFYQxJLYhEo3hXsXuEHllrs1OG7UCpPmv+nKkMXAXneVlhD
K3fp2D2ekTX8oergM7aCP1t0PGXHB4INrR2lcM8Q/BuyyitD0xaMSNjmtJvGiztX
neKl0/v158MoTvXGO9FWag7EYPa0jBqOiEOVMQRriSjCDqHJggeWogO02UrNc8Dq
5cgDCBYFFwWahm7Q5mzLwaQmfxthfG1iIZqFMm+daHyKP9UHjIKD0Wfz6FuMzKFV
EjmiieVj+h/svfgKcQIqP9eaPGv5eIjCuX5/MTv6yCIzNK52exDmccqCNGJ9qB0N
iJwjM3wHxLPkFLlHJ36fjabfdZjv6PQUKLmLHQ5XeEJFmDdCqA3ancv1OrK9+jao
2/odOlaoNrIGsS5JrPTgnVAhy18KwPEGf74exZbly+SFsjxYFkQCTcML/XOpa6vm
vzOEr1Wq+a9h0rPVzFpBHYw+nJCVcL9nlQ0Mqp0dXDA0BaNB0S5Ev1Ym2hSpfc1Q
Dgcy0QJJy8FWJfH6qp563yWJbC5EgeciCVAUQJMaU/K+N13h2OmltSd89vu3bXCD
VZ5khQdY/IupNlV+wIHyP8T0lEmuhHfgvjqwE3Onl9whzNPIYdR89Nwf6nC+TrfP
XgbYybL21W4VmaoGi64vcuSDqtuYaKwuhOzIlJx5kG6e64k4PSqLAiKQvCJFPxAb
/ABrBmdK+pfKDUgUYtYSLlhyKJFL7BEdy+ZtQhjx7Ngq43mmY16mvnRoLVYrbtzJ
tzjr2wnE4AmymsJfZRrNA/iVXb0vWRyVkrUe+P2QtcqQRbuPe/TM8/N7mBiI2yP1
210DxdAA8yChZy7wG4AdBd5Dus9drmL4d1j9EVEORy7lvQIrk1RF25hsPgS/6IRY
y0RDIKNfJPwMoHc0JWhWBphojb5DW6iwNJRJBLlvIODBNoLqWrQonKfKZdyw2yox
R5N/ZdA1WqoCFVWIKPvv4WUzlYGx7G1N9AkTqS+lkCCJkafejMyaDxUamIBGFCoz
Mx/WoKyifsKHP9qBEkx/Kqxy0JNpH3+5t2wx7dPM7N7AlfleY1fkRO53iIDLN4Jj
MymHgT6W4H5LuJH2saJly46ZVQYhPSaZJSYu7g1nAqFnnK0rx9o6zxVW0byPFyjV
oeQGv5wBM1RWCgnZcSdq0kdNv5hFCaYCHOEzrVv2Zsx2gQzcnX0f9w+b77vPWGe4
tzifg/vYkUQPUUJys85LUYhyGfegCA2beZPtqbdJn3WRC7b4W1zMgIBGJQ549jS6
E7RacQJklrNNizh/l4kWVSiQbEMgysUeuRy4PETvYcaOQYoY2Sg45V6FmHrno0a1
dBdzKi/vR/8s2+lnj3mVlKh3CZ3Le6lV5ppYA9HddliM7Bdy/xuFrsHhns4dNomJ
SMl7zvM4miTy1d5VHKMpM9fCAYC9Dytb+JUPIg6yAMLw0etayJ0FLbmJMIg2UYdF
1J47sw1ymYrdrl25gbttVAIqaFz8Qz8jhFzoiEaIBaMEAj3J0UcuCD5/HB04H6nk
FxI79+zdpg30A1h2cjySecVKNNiq/CP3HsA1pfFcyHlIgUZ+wKRK/QVdcF8ayEfZ
O7S6kmZCNS168FOBZGfx3OKolO0vUca+JLGSJS4g2FS9TLDepOLYMBBYfbxOOsQz
BuEb49Td+S2T9ONDsTblfW29QOOpc8+p2ylRRa1qKdGMjxKJd5vFmarHh6mH6IhH
8fDpXvrbgy9k/OqbSeeeuUhKeJIslxGBVw+JkMVD6EKNVbs02NVPnoyKrz2S8ZGB
VPvI/EMrGdyTt5BdXYbuSl9Aw8BnjFb1oqQ/P+Cs2XJsUASsgL/hXubHAHfIQV/S
bzWNSYwcECf7ZDpEJ83wxIR3kks/nQUb7K4N1LfXDZX4ZHsGuekpesCY/KOFNZnA
mVfLnA99K4xcsAf59cFZO3TEJmGoEeT5UWDfsQDL3uBdVlTgQGQ+hah2S80AMj+y
n4Xmg7Bo0f80yVfDRaIkYKfkgSY1ZeMoQ6RACIdAKdtXhvFXJJAohhzKthxH0tmL
Glesjr3942t0DTXG6o6ENUtLhlHUfbmaXw7AFgYRpTYKZSi0EPM2TvYfb9Phq54o
oCI2C0aDHcfOR/qLn2x4MuwsnrFTDguBcEKxQtz8X2KkMFwxcgODXvL4ZHKE3neg
n/G7e9aBws1AFKMIPIYsyqy2j0MP2XyXBlHbblUzSRNYaYT4KXVBACSnLFDqP5iM
igVAfDs4MS7CurEGSqGYjO6+yP7b3vcXCi6HeC5DN21XKiHTJr4i+uOsfXDf4Pjy
03O1Kh5m+vGHHwtUiu92lCdwQ+OCFqq/qttx+zj7sZD7J2u1BqFJ3A9YRdohvbn9
eWTTtFzng2HzJ9pVT5w1j3jrKY3hftqzyj24MFw5uQ76AkojEJlRx1j4QyWpD8Bn
y71lVewL9zwI1B/RUT4ZQr8YXcGhF2OU0mNvk5Vo+xPbRNVEW/Klc55D3y5h9/YR
kqayCm1sMhZlbcAVdWBCO6eAO4BNfFRQ0IBzFsKOKydpKD797Ke1DokUQqFnYYRI
dgceNd4pfrMRSglfJEwPbFv3qUr9I2Rs6Q3GJEQWyjH34eRi2JV2hJzDQRYH4BRc
L1ycdYNOKD+0pVl6/758fjWrtecmWa1KxQCk6M1aJj1lyeQO5nKh7H6jVDLprwsv
zwoTQNH5m5S8mQnIUbtdnMkCDX7r7egeCRTpbD81YiK/H50Ta+fYOiAw7TCWB7Wy
xYKh5wCHfhi/VqFwi9Xx4gPVJkzGX1dNktI3OUZidfwBBvua18MYIxWTomkC+I46
4yCvVctziv1iC9LecY5Pqg3OJdEfQjWYVFSGUSAGNQ/M9z5P3udhil4y1dCVBtD/
a9F+raj7bWJorOxudb+KZ4LtIV+utXb+tI/haOyo9lQtGqZ6ptqT7rceH8r8WHuY
Lsn2jAMardeLeHmDk/vHLZPbNqwrig2Pmx9son3tgRqyOSzRb4HlZMpRH4qJ01sc
YZpT1O4kT9dJ88oieOTIQVMoArMH9guiKFUb4BBQN88Z79rZVQ4S3ho0HmiG6PmN
2DTBBx7uqlOcCktP+i70DpXiYr03QRGbjwW1Wws69baEjpqZ5rQxhjmo5JTPdSw2
QNkHGQ+zmNsD3wldhSmCcgyRfDvXZJB7lrLI9yRZpRlKSo5VN4QnHTw9XyNirVzd
DKqhDk4DyC7v81TlRbnZEs/qXAFFnnTO6uQPKgE49GmRR6G7VMnh+bYgqIGYw8nH
UJSHcc7QQB7F7gsZ5LwgJT8PQo57uilePFrvcr+eZgQ0gDvbl/7KR7z4pEr20q81
bb5Dzp1kTJsAXr4pc+fLLoNAcMrLtwKbV+JUGwd2Hr/raJC+w2LCB/7dRGpMKPzn
FjETsFr6oz50YoA05/kCdgaNnqYv/e6j48QjZ2YX0Ut0MNMG85BHLukuYKceCW2P
Nsj6wL2vac0oGaCOwY4foQtUhWNK31bxv6D47BbZLX2YLl202gCqKVq59jZCEBzU
lpP3ovKdrO9Y5/niLy3qjRqANDUA+mZnUWoZ3YwLaHrzSZcQEwfpdkX8dumIi0q2
5P4ahgrqUdI/0VPkFvYWLp71VWgQmGbgHOEfsWh7M3vItTP44rdhP03YYGUn0/Yx
9AXaH3ol3VXk+rbaI8GPakZai7BCsd1bsFowZ+0SjUUnJvDgSZdevawwx13F7lzk
dvzsPOH5BGkprYBo8/RjISCKFwkHMpbhjkiN8rZeWwy/j+1NZZBgL2TThHorvfQ+
gklOT1lNfn0qO7KjlDbiXaRyD4FHRtFy2MpNDBUoxrGUwx2SEEKU6fWEnE+clZsX
tTG+Syywgi0jK8IlsMybPNudVgwYlrXod7jYTfHxBQBsbl52OMIxFFRZx5zMaOHX
5voWmcXDMI8E6P059UnWscKiq2cLHqsBEwl66QXKq/VraGNzzZmjwzUdfEaqMxJS
K2fAWRxsdrb0d6hOzrteAa6sBaIoR+b2PryxBwfq4Ijsxi+p7QGO5mEnQklF/PIQ
MzW6qpbJRL7xKkDimJOYqJVMAbSIHPnwzW+dCVCNSB21bA0Pgzya3ZOyWzjyc1aN
U4/WRsB58T8ymoDKS3FGeFKExD2UXQDdYKUQtQenagTDb2WNWpLGxWWlcRHtrCsf
5V/ovcWpwQLv0OTrLjxhVvtcSTjHhV0oxBgbbN45Qg81NJe19Mwg5wmSnDNYCMIT
vS2b5bg8oNPwfSy+285Q0WWwBz0InG1Ty65liEfJBV4l2GimjxryhV8fw3mXvbLa
X+JfiOjqS/KOK1WBx3krkBenkUsqKsBFhbQ0Du4GS3LNn3O1ri4wa16odtw35FYX
zOudNOJW24LDkgBxldZjyx29rH1W7pYZrIU8VzwoHfC8/U+Z6X2kn52QSjkUVGGT
aNKK/7deAR/dQkgSJeVMW6MBy2y5FwiGXhFOvPjX1MKUvAN6W7xHeYy+Y6wKbdjP
fwNg/V+6HvNuv90CIB45cQb/6gzkAJNUuN4x9mFWErLUHgR+tKcJNe2g9B/s8425
rVN9QPaQYyiwo0z0mZHEosPT9biNGAGlb3Nx+dWetIgEtHWvzzPN/lXTR9x6GeO7
/OoJjIF7sq5D/X2WurJCxECHDB2TWttYTZcf7c1cRY0eXAqwZyCR7z0q2KlMriO6
cc1v8tJV6I1sjr4jzUeiSIZEKEq3b1EQTNGZ68kG8XY+TMiKd9H/PFVIdq6Y1Z7E
RhLLiuNqj3KeDxr53uEMzE9+RLnWim0ObUzRIsjqposTPW3Aj+e2p1NwthHtuvzQ
JLxu6P9q2+8Vd6uXQEU2fus1i3r1SDCFvX7f5jJWKKF8K/L9MEk84CBjThiOEQd3
CWwR4f715Ddjj5tGUNDTnQbppsf0rhY0ZiFEHY9sded42Gvs9Cx7c63QZ0BJ91EI
ZURKX6MwOPRXHKF0mWbgmQhbhEjh9o54ge7t23w5Gx1URiSQlt4eTBuxve0m7zEg
qaW0CI91kZd3tVVlQr3L5E1epg0HeQXRzw036XVMlKqdycTLNipb7iEnMEZbN9wB
jp96PllJXLaZ+S8hS10QXcQxL7Rs2ivtorWfxwoGFcXNSA5n9aNs3Wbf/tsYbdE+
TrepRYvswWgtTn9Thzh/7YghqMbHCbKr8NOlt3/Hr7pCXMltdmUqYbsgHkEk3i5Q
azQ/J775MEjeRK96JmrCQHi5DdmVkHIMs9zwQZDbQE9+AGN9lCS5wkTcr6Hbfg6b
dFeZzBkCdbZ2XggavQNmmOr9axeESjMaZKzEO9TA6YSr9mPA+HUc37BIJ+GDY0v7
ZuxWc6M6QfvpFuxh24OoBWz09yvSIjt84Z93DJgdV8cwdhO3Cr/zGIh/3lQmmBeM
lL/qoGpLYIC4+9C+++7XyyewJ4f9/QFwxXD7v6+duis3Cxegku8gB/SL4jGGhnY+
SGDjOTexe3QTd0Mj9s1z8Btk8DM9ZKUFx6W4qtvTJbg6iy7UHf9XLvzsGTg/t4AC
3yKf3KODVYmZ14+v+qMOCq3zZ3BfkwIAKPM9bm1ft2NpgfBwbcdJqOzoQQ+WIbtK
a/4c2ZQE3pAPdxIkaqg4JNSVCYubIEj79OeJhCSsyfPlgRoA7/xSAx1YbAmQetG0
KK+3PudL0HxRV2RiOFXin0GR7CJTSeMgCOLuddmQE8l4efV1ucin2ONtjp3aiEbc
c5JlsaoTCi1c8odRaU89e/rHBBMW66EnU0gH0loXOExOavJb8AmnP7wiLJUhyYbh
pKpYO3Qy+yftTKkUdV/0H0loqweWOT07iT9qqKqTdnH/jWySy+VWhSzTdt467jHP
CD9NMSqY9c9llcHB47k+OlEpQR3wUmije3MCPnFYgX42+j1DmMwi+HdOgn4LskNf
OLeVr50/6/msvoPF7pKYxlIt2w1h34bVBFRcTFssJ/HbRlbuvNh/fYBJaTQlKTSU
W+CFnj3GimqiAa7nyqOTL9FA1ZyJLalOTIJAUE1mfGMN6Ma79HZN47NR1a4Xj4TM
4PJdMUbOzmAVK7/r6bGGjM/LtfvOoWuobfeU0YTf5z3A/pQ3jLjmuteSXNW1OlRT
UcB0PA2sKTzHXEtx/K9rm3vjvAfJ69P69UIg8Hsk5dZ8CL+bVbF4ck48knL/xHjw
zUXWUu9ac8r36fESWMe6+hyM8eQo4IbcGcElkx2Cmrcbtnhzfp13ZfX5kTRPcx9i
Zk8EJEzpHLvayBKHEZAk519aJ7h2khXZy+btPHxSHSoWp5BrShxaGgc/Px3mK/V1
1g2JqFb4uMwBBUjv+RlSu7SkdCxh/nCjJj/DMb+QHtnzEaQ6qBHJDVl2gfXbBeqC
W9rhLtq1jPKdtW1U8tqkKjgk7uxHNRrAPtH1uYR3wtYIUMlzMTBc6ilfMgRAx2WA
PjrOyqwOS56zpngQy+MBNphyCd1imZjaTlNaaAYvghbbCJUadpUt7XTUCUReLErs
nfP+f+Om4/xjjCFlOh0UfTFy5TIr5iXzoMOvSDgwCBa4aYRrS2yiOTr4VeGXtMS5
gts95DXKIJKueO4T1fJM41N2uXEE/0uFPQJ3aIP9LvbLEOFLERyLuKDjfu8EbiH/
Yax2H6pjbQuXD74QhEBqk9lqIwPMEwOAeLTmRWZ7pz7wup5ewoJSCOzsDH5jiLHI
IQk85pAPynnGSQFtoP6okSFUfNRzWOs9/1v2JXSduDi3Q9msdhWAfIIzJ5Lcdkb0
KgTOlw2qQ2ZX1kJh+3RwFFqMf+WXBfyNJ677GdlTVXj4N4QXwkwthB/kRkzvC68k
beIXDX8nfhjAvCjKApfGFWCn6zvJ0Vw7tHDk8wJ4t+5BVBtHEEM60HjAfUilVjds
h09QypIbWv5zdYhYGbMYbhksC9fdlLhXO7tcuacCjTW05VEePX2aOIaYa9pPoQWi
K9yYvv1a8WVOrOiF4VJgdf1mkUr7fj6PU9uv6Eqbg2yyjlDrKdeFhaSgtubCfFnQ
1Db8df/VlTNcPPBpGN8wyUFvG33shr98qGvj+2PevNS8DLO8o7Mms4FB6unbz2uN
/RF1KdTOF1Ib0/S8U+MXl5hUVCLykLy/yCtJ+5ieTsZau8dbk8SG8Sbl0+P1guU2
21vb3cEZiXiDWmTXyuvvdAhjJk6gJ70SdZWfGo55CxETDTDeuglUpY1Z7vpBkh2g
eTo9u/lw1m/aazJBzNnIXcuoLVKMf0wkqg95Uki+svxTIt9WbQRqFhwUO9IHKijW
La2coLp205WxRB7RSkXgU0q+EsJS7jEDV3Lg5s7OxPvy4WBv6cHTPvbo8xcDxMIS
AqgYlOBTXdbMBS8qsQJ2/E44Mq/e47ZutQzXDwGt7fYqhbkuEYCeHx9pNINUwxws
C4A7GRp7+RLn4veSQSKC6GKT5+QhDc+ex3W8Ew1nzZaaA69dCd6SILhoUD2i9Cxv
0SNuAgCBsCxqmHDTTeoS0esP4v8NUllUaVZv4+OqGpsjM5no9Qoz6f/w+OCR/F3y
J5lmixOp6XZdWG3h0zBqhsDkXjqldJhUY6Un5fmWDEdjcQa4EB1Hpgdza/01K19B
EOFyd9f3tpgpp7Dbw/0Xmml9aZBmx1DWNFosL5x1ZrHR9NvoJDznlTw+0ltw4eru
p7WWBJ/Ls4aWgE5leK9s0PArISqJqMUkTvOIekIp53q+QK8yutLunAe8rvyNNg9S
tG2RQywCs0dRnTYvUGZQrQOl6vJxvELyQ+q0SdGNTbvPKHnvsFMl2x+r8Z2pCusa
fPgJgC6KzotUYSL5xnQIjOx43ENGdV/tgozpyzw6icMt5JqbyMM0Lz6y6DAWkLN/
TULPQeQFDuC8kBRYwJdWDRtM4WuMbu0j5SJ/IHsumH7TtkT75Qbi7w3vBPsENNz/
7h2eqlV48NZO5Qvhfm8LVR2Y1WV+TRwcTV8gnJrSks1myHoinu6lxVfnhl6H+YZu
5r6R3BvDGSJ//SDPmECdnhjPffZBmU8NahWhx9R2fkIdA37VEEoJlUjrhP0FTOVa
4KZHkn7fa83G4lsjFExSLCpR6Epuc4r+zR3Kje1JKXnUcykmvoYEJZNFt27a9+82
i4eb10o9ZwNFDD54x137ufgFDv/ODXhh7mX6cX5uDB1f1E/iPRqqinjMTSPcTSsf
vJptKB2ACRtU0UcqA52tHSjwQQjrolejP5OJOnSu7J/IkX5WjPPSL0bHXv6gPyu3
9qtXb1rpgPYyWzwtJ8oaEWs7TJfxtIi1wC97b2QhpXQ5/GpiYnP0sOkfXV4IaijA
duKcPX27J3r8Suv8w8bmK22aYuYsOG5176Xqv0nSn4TOZiPlmzu2IGDc21kzdFNG
SmDEjk8VoKkFyrv3/mg6FveWksiSuNrHuUMnPknJm/lLlIAv9Ja3X9PuvMrVWF3q
bpNPOQgnGRLrZSZD2/QuO/k7y8VctXf+Rn4R49kzI7/Fs9jYNdJjIf4yxMUL+Cd1
3S57sxqovKnmoS/puCi5P4EOMCqXs2+CvbVqV9hGLRHdHOQUmBYu6e01YJ3NhTP6
d+ItuO7I64w0jsXB3Us8aYhL/jHvWrNjVacBKkMSTZV02TL4j85t9fcwVJj0HQ0Z
bY8PX5cLd9qbFtFtctvc/3OREyDOCOMqcUBgeVTCby1dVuPqeLRMUO6HX1LvOHK6
ldxHiSXnomtz0tkFysa4F5Fx/KQpxDB8b7oULj0ANurNgcHfzmFs2ToQ6UK9+dFH
r8qfCpOe6SOjHeqgqlnuxZ88j6+RuilSo2AnMGdGBmnXG0IWuY+vW/we2w7Av1aT
9L5YKXAgD80/CIB34jCA7HJAoKMzAN1/9+5BggChc8pfnKeDS8K7bCzouBqHptSb
cHQgkXUYvQpH7s1YB588Y71rq8SE6he99voeTJ9woxLpvSr7x6Y1Pu+b/uP+Sw3k
VT/qbf1qCZ4ixCDMr+a1FBJT41a5GWs6X3hhHFDEGZtGjb6thcpgf/m14O4VHi3a
x7AvYZVIf6Xkmu/EcprMe4LbU5xODYL1Yv2EVgBZ3RlrenPGaeEyOMXGKVpKqntR
ttT56B/cgThyCJu5mnRVsijBSYrVG+SyLnvlUiiMLCsK85XHAxMDFIdp3Cji3ylh
DLlBho1SyA0heURfiBQAL9y78hf0dHol5eNIELWzF4/HU91kw8ZSzLW1ihCk4zAD
LPEdij39Ujmf7zUofUgO3jxypNsjSiGkdcDefEoeBPxtKGh4LibdTtqy58swskYo
U5ForRKNrzi6npK3uBXjrlWbdjkuN92ycAmM2/gkTghX1qCW/FBQQfDNU4NN4twt
1LlTqIRa2d0Dl2Ms2j7i0epRzU1da51/VKPUrTAbIsIdOFRE5znKt9fxs5x2ouyU
o00M+aGFtuvCGjy3Lr4zpsFqGKOik2HWJDN53MKg1jCHvndZCJ6sWkmf/5BsUeSI
o+Mt2wmkNjOc9f6ZDvi2b6GYm3s98GAyKcw3lZnwR3JI0fRdA0FY62KSi8Nk0wq6
OODp87CWPl5XnLbn/6dctzSZor+BAQGH0+Jst/NjgbSJarrImkzeHmXxQ5Tkgkat
ejIrz0kQEl4cx4t7g5Z1JQxnQmER7A5DS0tI5fLqzNmMN/wVH8VZ5HFC9YIPViim
9qJvHZ7IFOj7lyKbOHGA9f8ltudmeigjD93dUIZpJ6e+eqHhUxUX/syg47viTIHf
ZjMkalMFgJfQxra95sQ3erzVMJb8PC7hB5R0Ds1cgG9qZ4VQQ53nRq79X9hTSsjb
3Zd3jfbEvuyfUoTFUd41MN75jEqbmkkoEpesDZTBFz4oAM1OBoIHyMDW0saRAWYa
5fBQbdAxg9NUxZibsLIN+nq0oXe17bV9uwN6WgHQlovOcndjRg8VZxPAe3AyOR08
YaPzssfRi7te691Xq2Qb/crZ+pV3BWUyzwzlimG5obWetGcIk5GAVEDG/nr1waV/
031/op5rs85MvfaswhypdQ01AdjzQJl+RIOgG1popWI+HmChOReGB2yr4iDzjtbu
Da3/NdOfSuMQSx0jfV+sQGc1uCutilFxsK7ok4g4gIXPdcjwhweRNJlLnmcErxDh
gRAxbrvRO8F04SM7IyB6QKlz/H3RzkMU6PtuFDnD2HOHbr2ZLuiiMSPFU/ZVbcRD
6DNUvlAbe1aJNGmPM6DVUJhglSLb6qszEI4JhE1lzdqihItEvbgMYFr5yo+/qNJz
qvfoxazX64B31Dv+UJW3LF0IWuKSJv7uNiua2LkZVmoM8ejzi11wzejODQFg1dGa
0c854q0AIlK18nPnrkMk/lWZxmxvYHrPTqg26WaIHW7lUrmi8ANbKs9tyi1x19Xf
rmOzEQ2lwkU1VRHe0+K5vdo5Txyy6RINI95xtPSLhNDBF4cYfFjJ0+qaKdWXW30G
wpi1FuQbPxzY3qmjuN2jvioksJwJLJx8or3HwP+4ob0VJuFcecuMetgP4TGAGYxO
VJPXIuv0+rh8ZzbtMpI7eBq3BHCK2OK0wzCBYC6TXVCxPfghoXL+0Ag5oIloAOQh
od0PXDemxKspV8M8wBUt0tgjsqbo2WA/AyiTJbZRn2pj2pPY45vfW8tAIu4s5Lq6
BDS2N09FuC6Q5rS4TjrcJljucDvsY/ZtXn7pf4yyQOoEr+FXpxwgMua7tvG7q2y6
HpvEkKiyWypsJ+phXVOKpWQUxKnQNOQaMQYiHZmYdQ/7jDxImJu9TsfOY64/P9n2
iL1ojQv+uRQ52EM7kuHCuFG5ocvgQgwUBlcD4Xz8Qfbk+oVQbQqs3298B3V9U/oc
HRq+f9ZHx0xP52waLiyKQL1EwsrfX0pFOEhngq7LMMRfQCcRZrD1W4OABmnKQAGw
G3Ii5zyzjYuZAeGbfFS779OW6rR8BEJZyauSmYN6jywQxhjistBT7D36sbjGkRjP
QKnsnu4ZCdHoRdHJ9lgcut8JTCCpf6B+hXvI8QnBhqDfLOr+ECN/zqS85eGhiDa5
U/lYtuSwi/+D9WHMMhl7ZBN2sjOsnVb2obBvhDWvFhngOqYRxH3KyKhju55m33lP
zZOvSsbg+l81nWnPBt6aFUEgJQMQANhcnuVhWL49RIDVAWycXq9d+YR9uhuwe2ZH
xDcY/gQVEsLBNN2JrQR9vp9+/IFIz00QJrulp0TTbNg/cGbgpX9ypunSKE70jbhp
uswxokSqbZKG4Sq0lAB+0lv44/rRn/4maagG+85bDB09CK7n+Elkgk7qBY5GkBUk
KuKWJRORn4GKl+gJH2Z0p6YhCoqJYDX7SaDEtagfLC8MQSBsTytwfF2R2a7QAb1+
D4ZXYbrERVOgsH8ktIbLAcxRgRgrsszAAx89UjoiFkEDPiiyEknZ4+T7EU+yVAFR
FIkfBWToON7eZeahnrKfNf18cajJ9lTaVALKcEh1mX69wOGdoSavKMqf1nKIeBs0
Z9/9kkZ28CpjvGWog5vK6MxcpK0tHNjBP//dtis63kdCZAqFSRFDRLyXR0T+3Mj9
o5RGCcQo4PyUHu8QqzffH7FsIPwx5cevNOYi8onGPPM1uz57ZKwANP0VPhS6odmR
CcRNdQkfvN3rVpPP5u50pi8xl0640RrWkJhuX36MUjGbz1xSExdQmTOx9YHz4sSc
ZgqAusoCK8Ge0oMsTuteJX025WlIZpLBIO+QEf7hATLf7a6npsAZGT8D8IGUAEJE
jDyNvKp5VoX+BifITGdz1but+ih/F9DBcaba3Uk6ANT6AZpxX+8Z6Q3BsGUax38x
w2X6KodSt02sRHiXQjfrId/D1PqgWdMB4l9XP+8pQryfkjnY8BD8cXIu9INMTUit
VGbw5o6W8ZXz/HGdXSnY44cyB705ynZhxR9/oJdWWHuLiYYIHDKB/XVlHd3FDfS9
JxwuwgdUE0cJKxJy7OQFMdYX95BXnIQDtP99ylZBGz+0BIMrACwYzrO5mclAaI/V
fzsEmyhhYeOCMiAjsRI6PIPPgSOqKmRnDnojj9MSOJEx9W+eijOxCAP3J87jd2uT
PxKynLOPLByeTeylwa01txXZP5UYjnEVwK/VS6UfzHeCRl0k5+oLh7RR/1OwELOX
kzaLJgel3J1KNNQqwaGU8WmCM6sf2ikZD9AE8xmDpzmDWGisKeznKClZJ4TIEFo8
X3q69xdbsvTCx3nupNmif/LocxhsVGV8LPPzAL+1UIvya5eAN4vQXX/KKNZx/A1E
mizYpOu67aHwuaQLSzlaoRMVCVSk8oEjTMSsGdVGNgZW2FNu4PH6paRgsT6lIfAV
L0ZwJGYbTIrj21etP78v1FBszy04odL8fmV7oSHGNAvhcBPELFHxESVSpq2qLPrQ
yRfUZs+5tzKSFDxFEWOrH9beT7VkPCRMwtuDUUW6M+9D5Qwc9NicmBvrmA5Lek+B
c3gD8xLvXB8riLjFCTQYNby5n1YU9Jey/tj6Mj4tHUbIbyVsdeZxNaKXHC6QJGVR
YCmGb2kcrG5dMFUgzIFvfsXn5mwjxurgWu/NM4qXWwl/i5++86RdcqcBzTE61c/k
wiDvlt9m4aBrUG5NGPyGZ0GhnLT8OGvPezF4ESdTlkw9p52dItc3gpoSzQFVJEy3
q8zTv2XMLI2jv7MgIIEkLB49mJyUYKHhIItaLhcZ8VEwbDtXGPoVgBlYtcsNLERp
Mcfixoq+P1mkVszB51BT7NnYOrHL6rk2yW6lxlhtUkgnjPr7rZLntM5uFXqsTFeg
aNjkqrq/xnzNvaU0WZIz7k/ErkA32QDaRQs0lDwVuHuhLl3K+xr5KBwygfY6MMp/
czSnOn3aNvL5fimA2uBSyk9WFpvl4CwGDE62DqloZEvGty0DrlmLJbHtmKp3Agbf
JEoEnj0exIaZ1/i7OnQ9goTgDgTSvvmlUzObXKioBjI20nDr09+27lncKpm4fTHr
sV2RF0gpEUqQDHsDBt3nz+GYMtjKzRWXynw3qn39p07vb5+lOSpshbxqd+ivStJO
oByDGfRgin5EiGEy4DoF4H8xcrwxYSU9O3vXgZ+v3Hw=
`pragma protect end_protected
