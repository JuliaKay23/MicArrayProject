// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
y+yLCjda/6XUzOH94G6dcOqCxY3oeL8EqebCBGDx4/My7riwm2Yy7uFJA/I1YpFOYa2qQlYtCQy4
RqkA4qkysOI0kfBrimL4Jr1UuzGk+N51Rw2qn8Hvo0izJc6A3MPbFPL03aVmAWIYUvWGfUSy5iNJ
ZSOCLgD3l2evNJ3Pq0I8tD3Mq93qIx4+eeXhKYpvkCvQ17F1H9qQVGv4Cs7y94OHsEBgZpnaJF9u
UyllWw9Rz+3pAPchxQVlnCI6SDahdGhyVdAkM7Iz0W0gG5031TKuVSI0kR7n83vlo/PcodpkiGio
tZlTR4/TJ54RU/XWFgwsJVB/SCumzzgn7kVZ3A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17280)
fFOm83XhLR8Ph/oJ7TFtzrrScaRdngUX5RsjCM1KpRPFmwSI3/TJ6NJKnll1wtoCWN9gcLDoYK74
QI2azOsfBGOyr3DjDzmEwu/Ay+CBdsdaRyjo5qb+87VJt9lGULbI7QtE6jxl0Sbhf7nM7eKhrA6r
oNdc7wEcSRCcZsd48Z/qoIzLDGIfBXwjkbrJnrMPqHwNSBvguMF59SdLejOo/HDLEl3T4eqhAB2J
+7QYV8FWvDfY/vQtF3TnHOGs4ht7tn7OYq3nZeGBcC3+SUqFciAI+7LhQlLQVR9jMMhTegWobyMj
Klkb3Lr+wiJhQHc+eSQ+I5I4gK/DnaCmJgNclTSd/TsPnk/0Jlh1ZdoBeJePmgdVCs9fx8mmVi1A
oTLUr30oPLCiuoyI7VsOSImzHfg6xZpTRWHJpuLWSTSNdu8mpxm/5qRIGSukdJcVtrXtirNKkdtB
zLdBVCGXw4X4ceilm8WdDGlId6N7y1bhMlwuZBYugbAiz8z4NYjDK58BlbwUEUhdif4ed1k05EU5
Ddl6UJl54lZbXu22Dh3tn2o/iE29t8L6q+0+7Molmr8WRV8KfyAisKKwMtBpm7A9sxsAqGOoV1rO
oBIFeOpfoST7JuzACiAKaNrAkb2NZrNLYLdAN5T3qXemAqAh5ud/Y/rHNtF2nsANE8HnjI44KG0L
mBgK36hqZldkhScIEC5W2RkVuW+Oc9xhH6tRCV7Rqqg01lhnPsfWY+q9pBFFo4WLIqW3t6nuDQdx
593OF0gwj8cX5ydYXJKYYy8nJHIB/Wkhdt4gtLWjE7Vykq8cvXaIQXLeAES8EvSVBhMrVzTZJe8u
N0tDEEHnKBVQVP7aks0tgkMs8sOJsrTwWIekUBSJeNGDTlRTA/7//SMmsZYxsBKVgxhTPJUh6BZB
UyIDXG1bvpCLUwDzI8yZqS6f7tDolOCH3Y33l9PewKLriBV5OVCdKYe7LA4/jtUKtMD9n3LQbvMu
FPCsMOtvqCixVpT2LvDBXDwHXFOZsxqSp6Ka7DmK/jG9A5ofPsyOxvmWJaxV30z7+QFQYIy5dEQi
w8N+ROzx/tf/qHoRb40fI4wSZCckX+cTDL/F7BBkqdv3OlcciIgUUOnMcjZbqG13eohViEjOI7w8
aQ+fW06O6V8kBekx1fMWUp/g75O7FYD3j8dpMoEORDEtFGipMwH09LNd0kJxkkfjHDzhgitcu8N6
DjqmV/ct/ONfex68eqv6d1hpeIuJJlD5Pnr23+WFFg56iWkoCa4aZdCffLqZ9I+DTtwMMz/AjMfi
zdRPa8Ki2rrWevQkhBvXSU4f2VQizWpWgToUNpo/UtYFpToJFdeCWMOQ3RSzzLi1htdmZRIkD3Iy
Fm0q+0hRhYCZKDXHuUfd9OJnRxWtVLoH7BTqoMPHrb7u5+zz/KoRTWwo4YoUYrD32XKS89uvhRDe
RmUnOSc43ogvaz2HzL3T/ybA4mVcmviJBVLhjKigDp3lD72vIpYvGRlmrwI+gD3AW6BRha25mifU
TGO5V9AvrT/D6Eigsw8BzX3jETqaugd5NWxaQCLPnfi5UwlOYK8MYUEHYeLB7emSLppICyGgBlvm
F3GWs3GXxNUWsVdJrNkDvQP8r5mtKFs1g4gBvDeVqxRh/TGMTjamuHvKpq0j9QsDzHQMzDXMm2sy
hXnUUfK9DL0oWqp5HpCEitnOt9leSGeYp3Ak1X4pDnviGsr/Jpv97oTySZrHtNY8xZy8zyrIY8Kz
aGXcI0Lx78k0zql6oStKx4XqZTu77GW0X90p6GCVododderdQRZFC5/wNUT2vCv5Cd065rfNmo7a
Gb6EaqJ7BO2sBSVmcEc+NYotx+TXN/qvmWPPJSRwAtcMcFTa/VzSPR8hhAjikGxAJxzecGNxSkTE
ifqlRa265m/pdb4z1XjRfE29JB4exffSzmZVXItobtu4VpPn7ic8Y10C8eyJlb6YCLu+/Pew8EcE
oZiJ2IVSU/2DaGhwLY1ggM5mYqv8xzCrX9U2XEeSRcQ8JajykEx6u6O/Xzkm1brRxXtntFseBYSE
UUT16iYNBkSxeS4Cvt36FsXDorsPvySx4+0Ufwaip2bWqnKNR1tlKMU5GAakbIG++g3hZUB3MsCC
p2zAnrARVR55sHMUpcYvgRAFgJmp3wNARX8ElCiYLpgWK0A48nN6jv+UTixSQs3f67KLsUF2SmTF
xE9fmGvD8+A8bPFnm7jp5Qu3qd1w8IJ2h+TF/LSQ+7Hv3/QRxmUURTEC38Al3dwX6tYPwUgLa2C7
cUBPqbXNMV/Ywliv6pT7spIsmETlV47ifzox+KFSmkAqxwqJ2Qd6kY8xDg/MfeDV1bcuK3Vz1tsc
gh9lqrd0QmUenaJd+/ve6T/VDyYATUbOsYapgdOFLPOHkX5m5pZxWCtckVSKuKN0MuJOr+N1dc1a
wM75kY4sWTwDaYx0uwqyLYgHSF8k81p0JDqtRWcdEkcK5D6pO/gdViqrysAy/ivLK0ZAhRMui6/E
tMmH+R1RkjGk1UM+9Tt9tpC6FMX0v2JdVjlcK8yns6YzWXpSnnSZSZoKmZJc+9gXy8LZkkzX1gUq
KIS7S4beevI8kPmYkm3NoODjtM+7moR/iuimBROOPK7SfGga1NryiChqVW5YLkObhuYncxDxV7wp
xZHAmJLqiYZo9xt/INOPF1QRbxm4AUwQBh1p5wcugpSiflGieHoTLNv6WLfU5oJK9Ry08FHdCMrs
G07pDyb9nnhmbdrJiCwvVKa7GiwHphNV99ZDgivtNYJXfBAybmFaGuteZl9HzZu0+kyxY9G+qTwT
Khp7WR7y8TjAU7MSCO+UCJvMCtlBprtk9nmBC/PtoXsMeiS/wBsqHZmyHsDAeFbs561kgAEs8eTB
kyv/hgexyPxjWhazGJD2N1UHHJp1LNZNIEzJzk3o5y7Kyq651FzP36iUBwIeFfZJ4p97Y4lyLniJ
gdr5Tazxf1yw3p0oVMOedW5sOfSO/TThVLQp7MM3DQJCHetm7ZcDDk4uYIrgms1odLnmgBhSqPiA
YF4W0HPbrxHDFLBfSnMI8RDausYUmQZSkw4+nJixkKOepj+ykRVZmRkACYR7yUltnMLaulazURdT
Wr9SgUMwUl/T7GMjJYv4vdNyhRuO6jQAycq/Igo+GlLVO/7VZFKWbTKTok0XuqDUwglYXOfpxFAm
yraRVMnENtFmr0UyriG+GOG1ejsPeS8YUjdZEjlmYvaD1S9VwDuDc5FmkdEjQ+mk6WO6cgP763Uj
4erYHlxhLWJsU1dEBr5rb+xXzj881D17ysgrMB8+HaK6xOGwHYzoxohyxhycLW2CLfG+FSdCNGOT
sc1tl4gU5/QaCdpQWtyiImUMZWcazpzhPLwVZXKLgg8T/uukHdxIbbDvx6g/FTCPBHxLQaRrP+D6
IpuW1WOyxunUck05p3WlcmZVmEwH8U1nMYryehDe6BN56Ktnc37a1BL4Hrp2z2eVoZjNOscxx3dC
fOsRzr5MbbCXjHqOttZNJ2Dj2a6wwFJQbmODmazy4rNXxXcXphgaL9ivmBYdE7mR21cVe6YauPN5
9qRnnoqnMbGjZ4TuzIUwKVYnGckGqRTPiFvpnmarzwCGB1fxTh1kNP1myJjv2KNphayJ9wmtDxT4
pcPfmp2BsMadBeA40tzx/3lW+Ur9LNEcZ+R35WdNGJC8oBdOy/MNMeC4SZxw25ghv+zMa8kY3fCA
bmygUP6gaIE47QDZO6EsspGpHl4DMX3+bfw10c/LsVbHlizfUuyA33K153s2YD3ev1mWVXpyorG4
om27+OiW/AmNaFMi+Pmvdu/1T6/+9kTP4rC4uv4yO2K9L7MD2OKhSqJewU7dib1sz4Kl9Ke/5i7+
cl/EtDqZOjCKehKW0HevjTQ4HGIULmU4PrvYtW/9awJwhs7ZRmHJyqQgUxRdnUUGjoARxUv2jVWv
3r+9pf86ldsGu00YmmX8a0bWpaMxxHcbSXyIPw9gLHWV5L4m0oYMlLB0ePM3wncQCUM2L6oHlW/g
aszAiBiIhGXuEMFF7yogQqPtSzjkFHe9o2h4ezsqvgzwvJfd3DDQp+HlcswT/DJdQkVBym763yqs
EeQPAwhecaXNM8orC5UTKxNMolzsIM8QVvr7cLMbfxGmC0loeroJHbbYOh760hXXstFhopin10Hq
PQAqJGOhNshKDvFaYFcQc2ehkeTlcdUaZTvpfY7QH+4D2r0Wjyh5r7KgHMYQ+UHzq1aRDDXk0hwb
tegdobTRJI1KsiUTe7kKAJOlxI6t6mzpLiXk7AiNmO4TxQl0kFJ7K1KG9W6swpHkclHxCnksoJja
ViCbOnzn8fiXj4C/AedA9SSI1jOguCWYYzhUWW6J8cdub3lzwN0M6mbA5RCGOEJeYt7z5odBj3kR
AgaPcE6DTIgyF/XBR6GtgJqzZCU9dUG02o7CCpQEZ7a0yhwXiJbtyDSEZw7HQzDSABc82d3okfa7
UJK4fTS25+aYLOBEuH9jkzv0ySjIX8jFulEMpa1ytex+Ye0LsMVQCKnC+k/B36p11d21WoImPoX6
kzp6vxKWYp4T8lDkMVbBimaFsJQei04Dn+0U0sA+r4rS0zlRbV0LV0cD3F/sf/IOp+s3Iuq9+s46
CgfNbzX/6sUCYR5UaxWPTd55x3ClqGe1dEclCpDLhrYL11JwK8Fks3IRp9XDX1wXJUD5dhwn6Med
28nY7HbtbHbWquEWklnCmLohIpIJs2umTz1dkgjlq6sj9gnR4tSykZBQgPoHpsJXkugtvWNorbDE
EvTXv4XDJny0auZkKRMAk6x2ApdXmGOh6FQn8oOg1EihTSvnyABw83Pxjb/satUXezMi23nMUDk7
ou7nz940i/ddOMqbppQ4H9eCNP3P7VfWVfIV4/7l/Gjqdv/hjhnMGJ0qTIZfn9X0TPzmLKGiPM2Z
fLA9y11iGIAerq5KNAnJ0VwvuAb1FDK9Ou5jQ1uL3Hi+iYFqWHWW02zmsP6HlgoC5UUF1xQuWx74
LE84SWK5+yIRx2SdIeuPpEfROc0nw7LWjGEi7hyW7qa+Gaevus/CMXQ0BL9xv8c3ay4fIXcMS5iI
ULxaKqm64lbi3R/NZD+SIrEJba+mrfVdjnTGQ5B/ik9j1x8/rYoIcBrfGfCcC9IVM9EfslCo3OG+
d6vpRAiPcvqZlEqRSzA1FRqhPScytfIDxWxupq4IGtOdUeSnq6Bk8mckrvH4Cnv5LCUPmAqwv66C
zibWK+Hn28YhBw/qWCcWXjoHzyUOk0UEmg1aI3aygOSFB3OqpJ5j7DbcFRCAOnjhNcw2m/azpSm3
zZS+qA7iiYW2xKNklvvOCDcviQdl67GoCIW2mqSU5OsOM60MGz57ampz/IxPwLPPvcCoFoYy4Nug
9AaP01QyHdSCXMxbz9sngYEOLmMpK6dT1oK4ISlycz4/mijZzhXw3jKYsR5YwGl+VCnlf5CvSJif
NSmtZJft2dbLgVm6/SmkrO5srEjuwlxEwOlRlkEL90R4IEW8VQV92p7/ub/ljHfU/Gk8/Xn7hjXU
4/QM6lIQj/56o/nvOaRYuC+k/ty4TMuPYszXCKSgt49oFpOkqnAAyPAhpBBf5b876F4RzINljt4W
l+8ySsjV9lnljZLWSCoMz0t4luqDHWlC+xAUO5qlTxYRfGRB0VOU5Woiczfyt4D1TxQKdihNB9IV
XxoYSu36tS5bvzZYuFmgn7dlguzg1BuY+fu33azWA6ogyzbEum8L6wyqQ+aAaiGuk1KdptYHxArC
Wo8VzXc732zcgWUl1j1nxudpTJhfgv7M14V4VA1DNDwhKt4esOLhkka+mlJ+41KB7YlHrpaUz27h
Yt0+AWnuq0XrtUQROIsHwdNeVKfU8/hhC7V7rj5FuPejQMC5LbAjVWCvBGa9iCdW5TyHuaDJvPbr
BpfdwEzOTYZ54iQHpnmhU+zq0FCHIqPi/mSVnL5BT1MW4ObzSI1JOXyLAqNDdrK5ZQd+5eKobbDv
28h5nbqvcF9kiLSvoTi8Q51H8ZQfNuYiu2RkRDxGyPFcdPoYo3eksroWnkIgUCZo6/hEPQivZTGL
jjKfoanEuP9CeOigmg8ayonD953ZQWyKUZqgxGoXAl4sPYDZjhLAVYEuIr9plbRcGcUYe4+cnE4o
3WsT23ijtgpx4f9kI3jiwd3HKCGjSmMtQcVFhsAO0j8Pjdt2BHzda+M7qrrSWQkXSuQP8cus/P1n
qwDD2kboeG3v6X2MLKLPfwonEizrmweNXkJ5KguTtaM5sUPy25tmQgx86BQDUnwqjhO1YVbSeJbU
p6RH7BmygFzr/Mr+NSENsqUO0RSF0yvw36kxtW1kUtmTeU33wJpWDKr6pytaT8j9K+x/Hs+LBbfW
9jXPgZoUCFifd0ZoReH8SUIh/hjBvMRUPAu8qoU5x/z4D7+mqrATP4IFQbDjieT4bVmrEXJKPHG9
JcvkynR8rHlWHN5trtIzlZgGtUYZAzadTCTWMTqDd2jKsySGQP4Rp818y1D+FTLUvvivsiqKEnQX
1Jqujq1TNn8EkiFFf3H6TJLzrMFXt1mx6JeGluoEzARTkW+3NAnv1Kd9XKkucEekfaHiTiSj6HHg
U53TVayA+D/sMuJ/reTA4qeLkIpcWEgP2zz6Q+cfKQH2sO9NDgYilwwDqdKrXug2r5LpgLBkUCJR
DRvpn8e7xreL0n2n9Pg8tuYisNK8kjs8tJ3/Ov5nQyxV8sShulICirFnWpn/kHhjijQK+U8qOTnW
VMg0fqWVipa9Hsg0oq5bZqFp1reshnjHxNH5YnJS/UrseLFdfxPjt32+X7CG3HwNDrNhbmOGUo9F
T14DPbN3dOBWLWhus/AQ7wAdLxQWUnJsInSkYAyFyfErJIIHHEj5JYftgMUgZ37Ct+B2F4jRnUNW
Nr21K38DWwOV15tluyo0UE6/R9ZRHpnePeinDHp85qbPGY1R27GCue/EtgcZtDsXTH9f9bpHcEtg
3zeERLW+PPS3aFV9d0jOTOAA8efWqaJwIA6gMETOO3ggOpD978+sud3Nnzh+20Xc+bIfrzkIJdbg
3Yn6dUVfZ2hlP7FdhZj9NUQFu/Fgmds5BtpvHXh0BzZaluV1o0xiXdEgwoxEK7LTxpmQh0i6QoxK
0vcBGp2EMUAe9P0SUfsuzrUkpsJsxG7GV4EPK9Hp323qeJQVQHvB5YdoExI3Nh8xSjqPODG76Uq9
ueaegtRzxWfPOYSJagy72xlJspJVeP4067iDjS5/iaD6wx3y1tiQksJUD16is9918mLx6+tUk3l1
wx/1wi4I4R7ZI/Db8+FQrMxkYTLh7lzbFSnwodIalfnPr0KBK+pbJ4oWVwqhahAYDwMOwHdVoRPt
aBzN8sU8Z8MfNfw9pR9aSgj88m1LN+yW4ZxViq8WRlgGQf6zgJne1nrbvJlcnbq7JphSiCp0/N1a
EYIEZN51DkV25GdNnZ2nIK41UK8ed4bJwKyUuj85rSmiDwpdJlhrsexZqmYRJBRkczALURXedztS
pyQXm1GX1zcJZMogc7yB3V6O4TqycOXEdJxU5fjLbNAfB3cIbWOPts7jFPNvk7flRPaHg0ZjESXW
PPVDpcTeXDQZHnrk10Cy4IAMfVEYfB7zfflGMhAzYVUB/JjsxQmoU+33vF2wp2g0aL8NgN9y+ph0
ujgEzkItnYhtZ1a+Syr0JRK5QrUQxFgJCSkS7VkP2zAVEyzhOpID9BD0mdie5tJY9fJuSbmPA5Vq
st00aWiieiTPUdnNOEmZVGqi0o6F81p4DsWcMdreqp+E2OEuceZe/c95eoQi8WvPLBhqdeLKuMNL
J+Dt0gsla8CRA3vQUJsZl0DGPJWsWbYcNxJ05NGdff9KklJPWTvEZOHo9lSEyGk1Fb/54OhD1bgg
lxjf7JjF27k8KrURUYdZjNo6BqvU0K6jxe3IuxCyXnyjozHSjQYfS3fTth3NL1DBlAh+WFH2Tfbk
i2pL+WD0NB8C1u1GNH1i8TUQy+jvkVYM8PfRwUHTOqK/P5nqGvIILu5Q3zcPThyqGu+aDXPaWoop
TLWG+UMkeb/TEs2jb8Ym6JB7ZiQf2Uo8lGC645jE4WHn5WvdT2N4pG9UMghUUoMbMN2lZt7s5pL4
FvgmgSvwEWB8b6hXwcK8elT5o+adDc0lOunnR4gMLnKffiAnuMvKIkEWL6KJLTwnkMlJFuPF+65V
x3bSfGGCxuHHI9v82+RuHKY2MfuFMsb2+Hcc26zJKxjXBpWsoO0j9X4WvSinAeGSiZqoITEDwCGG
xQsmUIQ5TD/n6AOfOB/BTmWB5qNN6DvAZGSnCw8YXXj6gwwX/WstEcfodt1PRcJ/KSGxJYk16Tt8
USEcCqjGEC+XLQZv7We7MStg/xJKhuSpwMsiiXVuexbwdZnWGh6mLnC2algaN6Ffyukp2ohQZ2sa
j7cjtCIhfzsJNe23K5hvk8x8+VBsUcZpZY2WE1vj/dRXECM12pdbUsSd2dyycSt4peMCdpAWPPG9
MKPg8rLObVnCtm5TQ1Qx4sgR4S0P1nU1s3lT+RkDopkMC9QiU6V19Kx/+0IrxeIHfzGHYlMCb6JQ
7Rag4aIj8dQSyIrNf/Setxv2Jb0YH4NI3wmEPRdyWpCojKZ1u/iRt27xOrFK8zcY6DZWxA+YNFOk
kYFR0GkXaodroLddABhM/9DyPUo9WRwRjPWZ77sfAm/bfaT+eszJtVQWvXqxZtGqMAT+YYkmYz/1
hhnnw1pfPhmHgtf0JTY5Xxip8f2VCvmShadCOT8NSPzg9hLbox2oO56wsNoDMkGoqRLhfQh+dZ2R
NB9UQCJHcmKdEqjZs9MgI/41udyuJhXO973I9g8RUbpV5V86XWApvGtBmUzX0/rdbS1Rq7avVfTZ
pcoCjVtZ+uUE4j3bQLX6VeVsLQLpqFvLk3MjmK+uGqywmN7MrIO9j8lRFEyz1bI7J3ZGf0pT9atZ
A0zXLXroflVSPMuWT/sMrImPYJdWNTEBKvXLS/HAy8loFcr7E6iMWjomkMa/Gk6dbPf6dKdio22I
2txy95lwQ6Zq5pZeC10l4IFgoeBT8TCWenrMhW0W4UQ/W8iGUJipEd34KEJ64l0lb44Y2wQ32k+v
No+YsI9fFdO42j/4NpbpiOOyudRWApR4wy5JK85iyLDyPDDuvSklgc806CDqTEWtCqER355eZTsS
w76wWUWq0/P2CesGrBA8u4z2z8qGXncjhfCYQ61zRlDQSGEmTTAP0VFChj7aAMg96qUJUXE3iBN3
8Cxv8EHpOv7Am7/QBjCkcWSvASo70BOZANaD7usczGmZBH6KI4dOaHvPhfy2lRJid1cm3peN6xNQ
9UMWDUR1nlhrX7eBdWRGFXLz7B37x8pVTzWx8jIk43/eaBV4l4MsfLD+mCLZtYYh70atwQ3AFfoE
v3wWdsY9kzo7KIQ0CZvjUDPILaCHF71m2H3Mp2UQzVhH2SamgIjXrM9FQtIFtuXE/KFonLsHAU32
WKEx2Aog/z4JG+TZkqObvrbqMN1llQR9o10YNXfQzXeTs7g22PYfobOeLdVfp6xb7/3Vqawxb/xT
8S6/JxFiqyYegBfFI+JWgfkz5/au4hEv01qtAxwVyWkRdmUiNcM0VZBR4bK6Fbl66g+H5dcX+YCg
EPT4CScC4JfG+HesL/ZzaAy9Jra/7FsCW3GWVJnD/8ofx2LhDURGZH/HAWq4qoeSG+27ngcwO1cI
0K7t3h9ccqs49InmhZx/HfVuqjbFkWOVjV/nF1dua/r9+54F8LCEM2EUEf5u43RO6YM6bRRU651B
PN24Qcu191BmhJOt0eh6PEYeFtb1C1tSOjC7TNmdqSVhYGJW4cP+3CSZEfMpiz4seolNB6dTfPvw
QxG5iajs4cKdSgkJ375dDowFLUNcyOQLHZg2TkgUdBwfQr+T/mjzkKKKAkMKVX81is+a4NSalZvs
DNEtzVRE+fbl5vOM5nrasoo1J+UL7Rw7JrkG+lSli8OyF0zYdBJ3EJkF0GUs3QpEYhDE7ZW2jflS
S3qGm3nFEzs1MWjBMyTu10oQ2fdtPGadt9kJjUmX50QYtx/39sOl3y9k429m1yB+cFFKfvE+kNni
IXcTIl5r8CY0QPXg24LVsK01mCLAyCD5TxktlZ/fv+bRO6iv+cQGE8jv3DZBAEeQlUFTz4QOyVic
rYD/CVnFW/z+c+WnWTqAGb98DDlD2Dym37g3jgOWmeL5zx3Y+Wsrriz0IVK8d/LMHOnfddBqQxqQ
32bdYVkyvfbRATpxxj3ox6larbY+QR2uK6uDENvMVm7kLrzl9VALP3ybgqThZxykaqELe3wodze/
sUQUHwUK4pQOkk1cMI5IDtN7v+8PB/NZ4SL8kzxbJvRP4Qb8iq7lzZFZFV6elTlte9VChXgbii7X
NeaBe+rGCeeY497Uq0afhV2PcXyxV2xyLDrEaWIIYbBX05qNbnzvkzNfU8mVlnYlnfyokj+hNuKv
4TzJDgWceDaHXbKuXGM1XigeNPvIXJsBkkRNyatszZrQxB7KaaNf/76WVbTdDZ55er4sBw7r8+mR
jFAxM44waBNbEJL1cqBLR5SpOIBDw29SSG0kS029zKvznDSoYreYEKft92QboiZd/bLc7oO7pcrp
8e9dGE6Sd//WQ1hMLSoZEIqXk1H/XFsFX6k3SUAF7kPmnwwnqv9DthHu3DK7x8jO0dJIRUv/l0T4
8Hd5uY8Uxh+YnlrbNTBlRY6ehRc7c1OuYmof76Q/maWLhsJlKyJO7E5DCVRSKmw3Lq40cq+BOTk2
WYdwNx8a9SN5QN62m2/LdjzSuR3RQE/L1QMGdr6Ch4cWzXJEEvuqF8U4N5pPNIU7KPoNxVifSM6u
JFFmqjPwFycgDtDv2v54vr/aUx3OAEG5KkuavA3bSUkLAh8tk2IU1wW2ywD0iOeKmJz12YRClnYF
EGW8Bu+LKNXB+BGQ50go4bJsUw6e8IySRwYlhYuei5T13hlWmcFWi8iPCQF3a9zXdYBKIYebuP/N
aeLg+rcjLMzQzDPhkEecu9ZN//xdREPcnaFDfS1/gjRaYaalD6lt6SvfZLskqDhly1+RvOzDQR0n
ixOqIXpQ+OvuGrL6kDKUKmI2sF295anasqJrnRbJ3YsrO0FgqJhRV9ERtZugWR1TdgVdtkbePZRP
Hvz37foEofHOV0O6aEIjzRIGAq6wViVwCKMDMVVa5QyDOPNX8D6DUyeCmheJKNpcZLiZPpOj0NzN
HnKU0bZPm8mDs3ceZdCuEZLksl4Wsz28WyTmySDSXASMj4fxSARRsehwm+t8cd3o0bGV6sE67l4X
X82Rhdl7wej+aRAvbTTiFWjeRCP5iXdC3mrdYbi2WBNDyKvpMmuTYpnQHoqXTUmM/rdW7vBP2iRy
/ryCyZ0oEdfsmsolWUnOHQeq2G/4+gdMJfgvXbRHge2LvC7pcy5vVWJvowL3v9meUVIUKzNE1gUj
noKuZVtVe3/ZNQ0U96kKyyZjOPK4RtqxE7RuGXy2WYRIrhIiSOuRR5r0mKmguinKiz5rvjkjFdXw
pREb/vxLzlXCktLxCa2iA+pElXpoYgcEeJ+Pjekucf+6TRbgvg0ykMHwEX34HQhOKOsAUQwVS1LE
xA/v5Yh6HjOTxD807ZqKxNGJzrxT6LrpV52S9S/7+EN38S20h6ANvTAIa4cKKwHkQRkm3Iq3p6K6
i3T7xIogrjl+HLgtIosFPhxggg3NLhblGQvRa84YpS256YkFgk78Nk4gh1txvVp9U3YmM4jMbWc2
eVvcIPEVhQYese20Mv2Xte21zbJTCEWFtMb+BFU8RYgdCRxEPUuQ8zuCyhi3Zd2DjDs8sSPDJdoa
J/offCXfYolf78RUe4EisQrM0eFnU+hUtaHMEgFSHWGI/taTymXqRoFtkdEH0IB7gtq/PPpO4/04
oQZSa6npGBx3I7j+isY6N4Sn+DUbObbBtkaAfO5REFSoGUoJ9rw9hH4030G4QTporRdPG6nKrb2u
cFDmfkZOb9EkmIMB9vU2XrnydntAZJnITb5JOY27kybkEoN7re5ZZDtiOJy3/zCryiaagg4serry
EeSWp3cbaRPTlxXLylkHcHH/uo/yNYDT3sJxbhNLXW1qLMr/aGeSFHZwNf8/2VYiSgDFnNNXA9rP
Upfp5Yjd20TuYApWESZbR8wAyfjv0gtp9/y7IspHbn+SyExNG5g5maC0af0v60pEAIMci3G+RVGY
YW0Y1J/Vy7exYNndxWodnAGzbhK+ZuMQwAxviBfTmmI6dcZ9YnSbW+W6klAcz4XwuJQWWp7MY1rh
nG1vu8zrOVgTpO/hIIpUzTKnB/hr2K+tNeQb66F34mt3ynPtznaH7/4+WieWEXGRgO93B658XSgN
pPOUuEMb8jhzcdOE9DxTWiIaH4j5RGhBYPu9k1OsK+m+CZAxP8OUuyqIKSpcr8LvUKC2zoDjkfc/
OXydnjHzErnxDF0kkl6aXcYN/2EbBXZigzI96IYzB2MJ7LAxsGXoJpRtiobnGRuI8b9Iu01trj8o
xTQknvkQHRPlW0kRDXGKvDV1y4adL3hZeYMbjqHCH9EGZx6RLM+Wb2oWDx962cjrbP7Em34qBepm
hW4TaZldLS43WYUpN5weJLU6LewHRHlzkgUTDE14SJ4D318xp8QcBvXGviqAWoS5TrraoDKB9m77
ub921I5UVbPn7KkI+uzMdEjEvw/l54BXKTOCB3zKBkOLmwKT9N4vpcaH3+bSMUp2Z4LsPevo31E1
btZhl0QxP6EW39h4oQTLyuPaChX1ZKPul9z0g4RebrXkWU4pyTQdaLBEJX0ScuofNYxz12Vfjwq4
WyYcVzZbGTvBCFUjfHF8riFPMkBXmYLuK7phA2WDOepf1l9WsArIlTWg1xhzlkZhEdvwS5GNxRUg
5RkJANepB1I2n67ljK/30iSt2tdo52ivlnOBdv2Br1XVilYc7lf9h9TQn/0lGO4C59fVTvgNmmdy
0mQso2OoxS0sJxO7passQGtuexApUx8Suu5tDmZO9RCoNzOGsqAlDGMYTnmENf+R/GCepAA3RqkG
E/0JAi4RIOBXXVPxB3be5iqUZ6FC7oqGZfpCA9Bqa35rSpthzNhKtD+TZ9u4KlGwP5aQEqqhreRW
uRZDKa1TtXtOlmvt74DiFVPzfAT0dEB93JKIiVW2l7XMb97TsqxzOz79XIAjwt4WUL2xQRVnXhNv
iqY+oGlCz+8eio+2V5G/ALNvQORLbmh6swqjExvO0W9TnXxbYBnsAtU0fK4tTYGD1Gamtm5c78qe
7ipTGGMA1EAVkzZLl8uPMsVz01lD31go0gVV0FJWTPgcZpBMxJulwWEjXJJsoz3WiGdhwhrzPyN1
qELvT9KxXXKyKpvemBzflbwjHUOiy+YfAOFQGUqTNevKpBx4luOXX9rVLfTDSgC16g/iKdQ6PJMG
cYg+4YqFjYpdcKr3tq1W//GVdf3gr1GfXovTGjSk1Jfj/Z6xWFfKIy3SxvSC233c/Bhwk4sVRoQ3
9KuEBIYVNfs/+/X+cb1rH9v+0F2wBzWl2eeE5SWN1Aq6towtNVuKEsPK69DDyKPIrCOU2pQqhzjH
JIhls72I2kgVjLO+1M9QxJsjS/ZAd6TwEG7VnL7OqKppGsAc1ug7BP4/1JIVzMbrkhmJtLeg38Fa
9Q+GMTduQOvRpCeJZ2SazRN2sTUYv6sAxvoVesFRsS4Qj36giB5A78DcznmdtxlpXmFMp/Va7ucX
SpGGhbu7XTFci6UHYzkUYGgwgLqenjj1oYbHzX3+hVeyr7Is6i2rcyojiA1ZmMA5FIKlJM3X9/bJ
ycGW+TtNe6SkG/LDs15BhqaTg2tpjZc/ShZMvyZS1VSdh41hBW03eqCP/aCYxJAhDIIJzAkS+0nW
+wTysuM6w4Z5X7O/ciLeWGLHdjGw8MTxeUrg78cqEiciwYVTAqJKAKj4d/pON63IX23ZQjBF+kzI
+/fYNEYIrrI87WnbDFxtAFCXabZ/TlQvWYq4vMu1WkYp8USW1PyyWXP1RKP8LmI5aHfAF8QdvFRz
ni46UHmPGRJh3MWVrsQYlWWdHf6XU9LSAIdhfBGfT45qCDObH6smps9sz6BwVUU/p31vG6LOqlsX
fxgyGVoXq+8vJQJtsBUXO/THrKhLJpRcV61V05fzEfr/LXweFwIeKgv4Nodl3oDbPp/g9sY/yJZk
maX5DQJweN/939CYdnfXmAeQqUkZwXHM1tNhWoI0mh9sUaJRDsuRcIwBp8Nz3Mry3zBfJHerEP/3
F2Jx49vIYbrBsd4IvOTuw1VckxuTCPP0tI/xRN3RYEXmbwMxmwNwkzxchhkpKVFJ2wJ6BklKrsd8
6VDDfPgT8M85WqmE+4xHWY4pM0JZCx4t3R4hNk1nkrnO55QKkw2utqRObrMWs8/AjoEn3uU5IcVU
3gK3do+KU4YYOXgKhTJq0dHGSw4B5YAmDcOPW3n397YDIhnxI19T47I9Yil4uVPX9O10ZP6EEzdn
UXiUbcqiunP6RUBcMS91HhNpjxhaqoaWKskZT/XUWRnaLCMuicEQmtt6+Cx07s3c+O82I/c8yweI
zRDzgihTCSoLB5x9bzOBtBGgRJgAgBZd7E6g1AEL4ZAIiuSaQnydaK9+M4O1NlEZkmk4PoQs3geq
hAIgotXknNjq3Cw3We6B7OUtrxoAiMZ8yjqgld94vWJeIVjEdPiD7Trn6VcYoEvlHMNqCvSu2bbB
dalnne6jllAQ2dud29aqToAykd6t5ceUMyPINkv/RM29mTjC0PD5gMgL6G3JKdaIEWnlui6hO3zz
OYEAM3bl0/0ESAgB0Oi9o0PzcG6H29OxSrya9PU3iiDgnKfLQaCga8gWx96R92MZr4Z1RFhEXbLC
O2Kst+gB2ilT+Zm4Hw+Kv8BhQyAype17C99oZETzS8PnfsQt2BlkaWVIn+9JHyLkCyjAjmNEdT2z
sKKF8fim72B7Ns5k9Rmoi4CrL2Rff/M6CDdN6ESJDVIeeR4EZ3NkKYqHC4dCGf1r9w8jaL/AoSBI
yZMu4/GOl68XoZed/OVABnvpkLHx/S74NepVgbGgP9Mhf8ngGEn7L9/qnLQJOJEIHnX2DLu5fmW2
xO6d775XQHIrsgcYOrDkhBs+440kYBE/BliGyMuH8+Xgs2c9o+7GryGEHbOj6ws6nV9iY/gsLzsp
3QVNAZNezbxl7COTKHPlOLqxrD4ox2BeduKD6TcsLC2tG3ufD1er4uG5d9wS4QlCiKI1eisQJzWw
Cl5wmR71vO9REkaoS7nUR8sMEhUmWph1Pne20nhhWJcpsz9/BZLDXyAzG+x57qJBMoXTH/ZhNxvU
/+PtYya2hbM++aJ3ImXMIRc5xgxgGUNqAZeNnJOKqtsxWd6UK/qPMTo9lz8qbHmDNBdu/XIVFM9g
uqJXq3CAgmFuILQDoDbH8S0BSKOs0pyGapn2Vg8HeDrBWC+s3hah/qHBy0rTUkFArDtgZunwhOrq
clQ9oRA3+g1KeFzP3hcHhgAOGCuFmtDydvHdmNje4fISTt86/N0fAtbldmQC1nDF4t+VhGjGvwpt
LFDOGIbNYAxZlu/ZCtm4TaWHUXVtOhRWM8iMRYnmZtg8llmXfunuasX76EzcVy6qdBrk6vvNHAh1
ZC1TTd67vptSc/fCz79X6UYqlGmHbnJ8tStqSIYoHBPWgx0neoOz+9drGM6vK8WyF+VHEZFoSv+k
Qh2CmLZYanVcB3b/wZlegti2tWngwGRkvYrBVvQtybdWloXCgNu8Lb5QLBpcnOgMyKi8x1vtp1x0
qfLM0b506oWd77+N5XVHy2VZ9fhFkzPzfrpd43pY2i1xGYvjl3yEs19hYnmUjMdfnxRIqVpzB/10
YLxOqlQXdWRVfcdbtEEXUy3IdnyTKdxz58R8OiqG10sAYrhD34dmX5IuWkJQLMdEobsq2hWu3bw5
ZBd3SOiqsonb1xzqEkoE+ZQ8O5gDCxUIRR/kD7TMEh8QEFISM2C5tTmYxAF7rSCNCNkOZ5x8h8zO
aZdQZGl2VQ7kFvi74hpufHvjGXTyRzSELwkWSdX0++SySNKyXYCvupoUldIrDIiE+clA+uJXMa66
YmIyQt8ETRVcl4OPEEpWHefNSsd0nOE+7iFprWKYN8stMuUZKjfgLaYRNRwwzZio0MKL/775gc9q
boKxvEQM2Jw6wZzBEgI3YRAgMQB2TN4QYFKjF4dWDhyLETLFREuDprJkViay13/0j5srah9l3mmu
zsGOkQNVRsD96QiBUhgAKtw47FWiKW3FAqjGJeZk2fimYPBHD83AkWw4SMRyqB4n0rANYLdZKERx
jeAT5qWWPWoQkrM/A/gb14sGLnT8LpXKNj4I259Z8TVCQtk/A1AonBoDjQYEST7dpbkbUopGIVe9
6YIHTfEPZo7uoI/5oNTg1tWgCcFIaYZ9dM9sqyKwsUYD4R6YIohyagBQP+zm3ju3Ot+RA7WBXFyE
wj1bVeaR+IvyCfw45/bQiRRAWRXuzpC2iNPlSzGqOiFUX7HZ7rT6F5MtBPDK/6MwAbaVDDpFydPS
C4ejF42vViMvNjDEfzXaHC/rA0x6oGC9OgiyqdZz8nD8SzQ6i9g3C9xz4iWtpxBwrt/IZ2bgtkr5
g4cv3pLzm37ae+KVQyukPDzTJ8EqwyWnc2NUTZB+YfaYZpmihENMmV2gJD68rywx7OJX99WrsDAl
9b7FiBiqmpVeP/+oBMZQx5LyZhVkLMSN3d/huw3l3r0gUXeZEtmRfLDYq2Z0adw+xArFcRMDTR/9
+Dx5b5QJElu7tISGUl1P9eU0vGCmLWjnVlZE4qUD8MUJ2weNjFOAHOdOKFu/W+Y46ZaDqa88nwD1
F2+p+5NtoNCmDtSM4BYc4LPI5pzRUciRQU2m9r4gZ2VTGwEeulgum8jhg0EjmLZ0ugC0Iz2o9SWD
Vy3ukK6skWwSlAqcbqQjmw59iMfLqcG4e8HcfYNcmiwQGZSoXgGvBwWcLVOAyoTR6EQuDmTfEFv0
ALbJcS1Byw6tpPOz7Ww9ONAV9Z4P7Y1uTFQpa1lxtjqA9s+d3ubP5dSQgpuZrFRa2T0SMFPRIDOr
2YooIj97SDiBxTavGUvJ92CxCO9XiC4yiPD7Gy4qGKT6U8/00ld4TysEmttPBn3C76q6FnEN1KvN
g6LyHc+XSQ2Un6cToZ34KUROfZmueq0Z2dyBFNzc0k3JPoJnQVmns8Svx7FWjFCrMD7s2p+ikNRV
dhWjP1UZKarG0V6Yj7DrsyPj5nCuBggSOAIREPXxHjx6NJ5xKy2dUW1UYUJdz/+2X3meHSqFucVW
b9U2yUhurVSgYY90IltyWpv566SVWwq3h2u5mppnVTkKnxJMZDW1VQ2p9kSsxvtcd4+j0PcoRTT9
DOwHbL17QgVVrNKCXGMkTTtJiC8rlIs3MI+zC9AVoTrpmCIj7hoYQ78mKA3MKOxEsvZ1X7BQqL+o
cqq1XJXrHzPlX+YLJNVq9dPsVSLKBAkM+MIIvf3mfy/ooeIJRMen82QsL0pmLgKZuC/Y9e6PmLmm
81882eIgRlzlSLchOPDHzECgNZAzi1BvmBDCysGt+nZbaa9ANrT/rApyLfu7KWM9Cf9OZk7hMSyk
wGJTA10n2aRIdyn95AjpLOfPyrC7RYvwEz7qN8VfJavhMdq5b+KJrkd5YPebQAqW1pYqiJlySzt6
7W6vCq/+bVrCREfBkqk7VG7w/kzfrO44/GEsLO4a8ASySHy2vepfknbS6gPC/sDTIGzX08uEoUDs
w03/tiQF2uYC9mhwqEuClGshWEIre5dcDSpZ5gxpLlDoPbZC/3/eselH5PQBEWB96pUdjU7YCnXo
tXDPyOCHwzI8/jR0vuoDruGhveBTi7/JdPKBcLChgp2s5bkN5F870yNxdu/Kh2TPcUjr4NQe3/El
2f4bNAZYcsHBoTzK2CEyHEjhzPaBR9BgXmKO7zkuS4KzFYYsG5h8lGTON51bV3g7ZpDytIi1EkK+
xpyT3Qv6ifSVPkcT1tmtsxSotxtDHOUMgE0D73aGay3uFlr9X7iKSu16XxXIBNrq3uS+ZZPXk9Nd
s6rZ4G9Bw0w0frGLguU5meJ0Lly92PY3mJjpt9v8nlP/gJM226s8VjFPvyJgo9ABaFxS+XeXE3b5
W0snDU59ahLrWLb6L8jmlxDEzQiQgKr7AMY1L4V3BK+AOKVoLb9vO3WSK1W7JLN5hHjkgao1GNJO
Qx+fqavfTslKjc5v9wExOAYfOkmh+Kg6IkpS9uKNI/FJO/QM3DSlqZFUnTgpEzJ30SlQXAcHW6nA
5ms6jSwjBeY4W4cjeNtz8+j1DOFiMn0486tiIbOpRmEPAGyF61qFIm1cTk7NQJIl0Hap/LnzjKlO
OHrtMVJUQSPs0eENMM1oPIBWC5MqNnhF6cXeULFd2ec7soV2nhSFy97BvsmFthSOjQvPh27XwfF8
0rkTcTnCg0CZeuVvIAbBsJILy5Jne49qtpDevRwGSJAjBQyBGBuTqflkgBQG20zviSLShD8FCMBU
IUtufAaUQf6HikFY01+rNRAbiQ/CA1+0rYBCY3wimJvhbszfX8+jkP87fC+g3ZVkTAWhQs0tRSl5
z7PWPWNbA1Vt2ii4DRcmkH4y/KVdcUT+kPGGoDFeT4ejLk3NsNUsOKZRvZeGkpc3ZFThrONoZNiq
lr8ZAq52rO35Bp7/waW995t7o9to+PBrxoaES+0DSaeApelp4nodf2GAaHMySNDedrjnbaRRywJV
FphCKYYrvxrCQoriYd0Kixm+ti2Yn2g6QudA/ts0RzC1DPzr+zR/pKskNjcDg/2+xrB+K3dwmhl2
GPzciAJAi1eYfajxiwsfu110WQXgaHyBd76OYqwvILhX1uMdaZuM+gS3n1OaD5yGfheYXEU79qD/
X/mf9gcQ9Rl0acBzaKke0GJMxx8XMWXg2ULFBlQwVUQi/hTFvnlrx/aJnAzjP8wWdjaVGuY6S6O7
wLY4RQfaJ7+C7SHZGrLGKGSpLAUk4l2W8NGdNtyYiLisg/KAi0uNK6oB547pDlY4ZfKd31i2I93e
FK3+uL6edJIgjDVA6QQUwgJxYFG91RtbiWIYICYBiyg6d237Xv8BF/4jfAp0tbztSjY3GTerrBcd
gbz0iY3U4yAAm1xG1UJJUxKlwhMwMq2NdO4s4yfJHd6WHxtC+Pl90HOE72ulrmqtCJdvo6OUYoms
xYv8YYiVW1cCP2FpPwss7VG8/jNPEuYvFsbjUODz0sUBZZccI730P/PnsUuLk/f+FiO2Gnb9khck
LkL9gwp56xfSfCkkqaoe2KMy0KuuYn09KBAXe6qZRyf0HydMHeKSsS7QOtwcQG169UF7Uu2vaWpf
ukeRk0tiXZOkfMtkIqV8myfBV1UnzIvRHy5oZzSL34xYIBKqLCEvpYBcuK6qMQ8Ek5TGjeY/ACgX
WsNNlOfiPQbGbHm80zpQX4tnx2z2WK+4MfWV329yf0g+2PFDYw+iJh33Ft1LS9uMV5IWiWNPsKAY
qL31jJGAHuBV+iv8VS8A9kee4IyOs7YXkwD/29e5/WGj07Kwn6VQF+PAcJsdFZJnuJjVKHrZliwR
gWckqJOmMAm6cuTbk/TsRNMw+5cPh5PkCXPRrlsMTZjVo+EcvfWsp5emxeU+xk/Q13gS8+xvq8zA
ox+CHAYKpCLDHLdrm+HDSE7GPC4c3A+pZ54lvwrt17er7zkwQOZ2MeKl3Bmd3MC7isXvolctH3tV
tFltUXHfVQ1tfuug7GmjLpjUfreR4phjdc+LbfM6Ot5ki1XcYNBUhLURTrQyOMbwTZyOwqtPBuUY
FbsPEVUmyprAX71ksVTFkNJFJVfS0lJwVjSPhdtLf61T05L6V1NoXCQ6hX7LH241CmiPGSgB1Apd
jn1UWnvk91neoXgjFyK4qbIRk4jVqN/9SzGwCGtOt96tie//S4t+nUDDj7GhRmNoeRwhUzlr3+XA
CviNh+sgOQAHJXoDTIfZeu8S/0Opi2yGojqavWfU9IpweGtpToNlDndktkGWVhLCqvkiQWyYpQQQ
XK+YsI08LxVAw8q8XmziKFjJ6cksCFghBqUiO2v0Vmm2/K2SQfHtOrrm4YH11STTQaeakPwL/TnN
8wtHk+QfWr5n5N4aTwCOno+KxBX5dSb2YDKc/mJmXjLGw/xe0Xb6TqvXupyfX6GzXgV7lmuv2zPc
3YzKWrI0op0MNG++aH2+xuKqSFN/z9T/vatjMbOOI6Z1a2arnyYD7J2gIwjGKmh2E8CLRWHoYit4
Pf7JXKFsV5xKmsr+7PO1DWqQsP6dVKSnueStz41N2aS5SdqBpHUZiurHpUbr2m6mfCnY1JMRMxKV
4xqNk6mzt7U09W/l3ltwXd9HTipTGV2YlGfo5M3N/SgpVZWnWrGAczmAzadqeUhdMY+pnjdA7iA3
PajOe5CX15LRAYd1QDxfMrB+tsumrMGcrHQkongvqtLG7cLMLnIZOtlbDWwQriW8u1M5n81qhLfD
OvUTkQ80sYKeCno6SdtlTUN57dZVHA0SA2SsGTfqskKnmOEO4Fj1l22p4zOMlJDukJN/YBPD5M1U
VQx6DLOGxZy1o0UJaF8lqa2vSr8wbkuN/cHb70TQVtQ9zPRnzfTsCIOz9L1d6pqB+2+rOK/3ixcc
nY9wnTGQJOhQIHPkHwntyMVsH9QdyC6lx8XtpCrSqRpidNf5gSM0tw8h7vQ4KUGT6EUw+ZNf4yGb
Tr+/3agfLJos4005nKoYDypTHDhqODNoq6Z3tqZ/JzKu8vNOth3FCTI1hBdNuIubmaUGE33hOdzd
xKL9zMc3cqYyrsk3bqDvOvT5joiIUfF0uHwA5LP9ApsPYYfZ9rbpQFB8gx5hVUa/XiErJRZN+XYa
TSJD+xLfU0FvKYAOtc5xLOqUU5oG5XXBK52ANb4x3PFY8j3KfWxMmad14pydl+jFCBXBcWty7Yp7
hy5eGcAwa4JMn3QALqfsCkZJPfzn7hFaWF9wDsczXWn6N/Nz7socsXEareJb0DzJwkxq/020HZk4
KM8i3VkY08PTPj3984hCDgVaKKoVfQN8Mw6qakfGfRdwjw710fWoiuRgVT/uJnMoX0VcYoSLSxA7
sUI+4NlGSeu5jsHw19ycAe4hTw52W0tMWgI7C5ABYeMB/udCy2+R7Qjx5jnqtGascRnuatLLch3g
usNn5wkZIUYaM2PRm1eqrJq+7gKmD0Gdlg4D7ick0j8S7coMiJfJAluNYhFXOc+xkQPRbGQgmSLk
de3mcF675n/drUrTY47qaU1R7fl4R0yiUhaGIOnqQckEkS2gbl1xPERTA22C0kEFR7LfWqq6wddA
NUympb7rdrJbE7iZPJIcT5OT9gKR5pZoOSUV/0dNH8boYNlPn0aS8eIbc3P0jhQs4VLhH/H86Ver
VaBvEKMBT7rOJOfuv4qOSG/Ey0XUOFQDkDtLQ+vCXJ3ZV6YalgTJQ/bFYmTO1eMpph8YIE+VZmKM
cQu8NxUO1CpnG3H2IqhHlOs4p7aEidUeVBpRz0M0ajUuBwdd/BLZNxwYOjj0lTZLt7HCL+a4T46w
DqVUR0qNd6JAz+TLfQYNF5eo5XBg1O/OVpHfFJdKC4OHi8IVdGX1nvPZIOYOhLBNDKgbdvVGgt1l
eAqg51LLclPOyCZYyZUZzGQSfXuqSK3WGvTl0RJjtXuID+MmprwOsSXKyLKLa4unyRkHRDMhfhgG
fEEJnARdB5O99lsbBtW5BxOiHBsXZ27tHzuzcP3u1DG2e/yQ5XEwKbMjTr1zwcc1u68PnmUOXPq8
H+PRr78FLwMiTVKiUx3V2tmZudx9dReY8EwzuNt6+XdGYsMJIMXOC4h3IgV+464aCJKtpiQtON/x
Z9pgTup3sbr+yLvbB19vrUb+do6iyiRZA8hFVRF4ths4AhZeIxYN/INUssMcqOVNuVbnF3SPxoqG
JbnhBynmwPdZVw4e2SD44Xr5qMJLhMTUOgSrqOT5JD4mq8/QR4ONlDT4ibUFLqtlJE3INKzUsQvj
UBFmXsk2+9OGyRVbe62hRjRYOKJAqhZNr8YK0HuFxj+AQKpmtlHZJ+Fj/thI9bKEbIDQuPNu/p4W
ACT1P57EPgCMJeoZgP8xI9d3kYz6SOhLm2rjpT1jVkBEOnqLiL1jsyFm6Dmbr3SXqqreNd/1lRLr
6y3KcPfzgQfWuQDLH2cJNWFPmIs9SQFgkl5HFKIpU5DrZhtT4gbDiuILR6+GMzrS3cWgvRGOEx7y
nBMc7Ub5ZUq5NXzZouNFrLFBfXRBg3sJAAuCAsvyFYCUfTTQFQb2+yS7G8OPXhnm9+8RxhJLZdHf
/sNthWWqssowWmajs0R0NC8Dxe9urywRb955W7pC69cI9koJ+V6f/k+udA9pCUQ4N3z4Vtn2mUt+
vYQph46QQuzaN1wEAOy6cTxeQQXIYo6Wqiocq4fFn84YaP5XjjZsnrGVfxnQXPet8zkaXJizVKTt
3vfwut821Po0aClzfXkQLt/xJPpjLg7GSmDakXdvGQJygAYDa3rENeIzbTCm0ceeXZx2PZ4+dW19
cv05NEIQy41sDwsBEs3cME9KNeOzkZ3/ML6rYLRtYBwj9EnDtQp47odGF+aUstO7c1v6GEoEzmbf
1o0Ji/CgFfjS1Lk6aHs9C08s3nN2ra5JhwARt39MhkxsAjzXaATkKdjj1A/yw6ImGEUcoxifDKhH
5KB2oczfzFUBOGb5zOX32IRlnsi6c1v9+0KJ2Qf74F2ZpAL5tRGJDU+yI2QAGvMOKABqPf0MHPB0
imQqiLcxQqBghZ8Av5YE5ntpOQ9/i1/5PZoPiz3Ci7i6nz0pk66tA78RTenBz1Giewu/o0mo42sD
lUH2Bg0AQPIEo2MOeA7e0nH1hs0w2gpV/QuAp9ePGgRQbHXIbYzBVJFg+seWH8CDKVL0WZppwpol
gOhGqiSubFkDSoW3KonPuVepn3ZcuSExcvLrnsKIpGvO2WDpw/xZgzVCbimV/7fH5zClApRDnbRN
F6T1epBYPcQ+
`pragma protect end_protected
