��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�GN�Џ	�U�1`����Ƽ����}%�^H�y��Vk�Y^mUG'���eRH�^7Lx�yq?�au���/t�'I��>Tfg����d�����>Ҳ�t����n�j��0�IM3��d}�v�w����{�Y5����eeJX�����r�iM�;Q�߁N�#~Q8'ý	釘u�1�S�Ź�7�tf-���� �¯�cZ�>A�/�"/�E��7c��%V���� ���!�P�<wKT��G^�P���#��v/#�8}�֤X񀐦/+P�����EȞ9�1y�6�����o�1�2�#��r�Kv����u�!�"�,Շ=s�b�O�Z	�&�-��.I<�s�ǲ6�:�M��&h�mk�5�,�^�5�	��L�#���f!�T5)��k�;$4#�&������Ԣ��E�1�N�c�'�iec��H1�6CVz"V�((����Y����	���gu	���_Ld�wl�ֶ�6q;����1r�N�B6�s��wœnI
t�0�Ø7����a��ǰ�˳�·Q{i��Xs)sjjT�֖5����d�TF�L����f�¹����c��(������o;[����$����s��ys���N��,lL�v������CvO�߃�z�F��i�c����i(SGmͯSª��7A��K��xp��=U�������/;nL7yT��:�?�R�|���G�r[}t�eg�X)���g�$��]���J��Mַ\���'&Y�aB��
�u�A�Ђ���c	�{�yœ@�}�>�+�EZ�!�Rǝ썄k(�@�t�hߪ�b{O�J���Aקg�u��b9�Tl�'Ȟ�x-z3��N�~z����[d��(tA��~$�d��)��b��=%�{�\+H�W���-�y7BB�ؓ���-�O�+�?$��p�tv��c�*��&;�Zl����p���	�<I)���fOp����xVvyw�c�Ve���H�Ũ�͖	������W�R��;P��S@�����2ɸ�%�Wv��gL��ZJ��P��K�#�D�@��]���D k�W�
����0������^�5kn��e�P��c�ie�Z���Đ	uI��=��E$Z����(��ة�gеPl^�5���v��5�t�F�g4�Z�����	oY�Xщ�
��u�^�s�8�x���[>."8w��E5|�J8*KO
�}��Ĳe(��zw��];�|'Ȓh���>�+�6��2X����z�!<k�a�86��!�+ ������b�p?�*����������o�xL-a:�ڀ|�[c����sW����L�
DT!��Xh�"
Q��>Y�ڪ:�c�[��ȣ�0�T(;A���u���糓�jYqQ���}������|����3"��x�=��i�Upl�W�t_�o���8QX���X�<һ�{��ga��9m�#��1�M�Z�z`���������B�'����n����{~����a����k��/��]�}�\f���� ����~-
�e]��u ��W]�zp�����/��Oa�-ѹ+T��p�D��Ҷp!���to�P�,�)8�޵�:��ifs���9dQ�-Gh�r�:����|I5e��Q�����@���i��4��]�H�f�4'�8K�d.��C�IF�޺:mR�צ���r�l#x�8[J����=��5_L�BZ�Էx&��80�X]�B��>������b�}s*�Où�<�o���i(�W����v���jn�����օ�N��q�y��D�O�O�L_6�8�c痺*b��mbt:���O�ns_�wI�}�A�x���6�W���l\��:�bt�7ad=� ���d0㗙3��Y�P�k�^����Жkt��[
����\��_��ho�h�N}av�IZ�ҵ�3��|O��<w~�����z9�k�3�E�b�P��=���'¤��O�*2���I�U���~5e� AeK�D{���J��}y"���No�\f�v�~�s��E>W��fĉ��{Z�PB=�����)*��U�Y:]�K�E�-ӳ�<.!sa/�aT�Uj8�=3�Ӽ�E^�.���0�2�G���D�ďsbU�)�"�z��AN�&t��(={-�P����ʭN�p�����J�CR�@�*Ey6/HR�
�@�o�)�Bw�g�0���s��H(X@��O���\/�F����s&i^�V�A?�ORN��˫o�N�)b���c{���t�ޒ��l�Z�{��;"y�J�!tj���X�F'��J�^�{c�w|�A6WG��֢�t #���^��6����-��?
=� �&��ƴx@Lu���@8S)��1���dQ+��m����n�} jj����s�j�R�,&Qe"���!����=���0�fŹg��zHS�9�@Gή�iɺ�#H̬����rg�fa���4��0����*2�w>l9G�r��������I�5@��`>=A�_z���*�+��b�O����3m*6R ���R�5E0P�p����.٦_:IVz�
0M�K��<t	<y������5�� vk�����)��*C���YW�zu?��FM�`����:��Z7h�L�b�!�l)D@��	Rt��U��w�@'�)9��e�����4���A��FP��hyX���7�|뻿ѼG��Q�Q&r�JTZa�T��"�GQL2�C	u��m��.m��-�|f]
���'~+_.�2����$�;L7�9�*=]������C�Q�tZ����谗��t;~q�۽/L��S��ӎ�o�6(���>�~3��+Z���9�+�wE}d_-�7o�#��t��A&ȎZ� �U��0�lX1����_g�l�t\�d�2b��%��L����=�^�g!�at�Ef�/�!G��㨞�]�-~ϲ���Q.���`�]8��g�G�$S�, 	#�,Y���ZD(\V�ђK�8+� �';t� ��Ձ��D�5w��c��Շ+��D�O�eF����O��≺�������OJ�������u�R��C��7����6�j��1�$7��8�(.Y:�{V�-��
���f��zSt�|LR_?�t�$�(�~�-�K�2�&�c ���R���Kwm)���/�	�o��:��Ūm�e/W^7-��6NA?b۾�$��~�&�>���W�ۙP�ުT��9��eL+����_�j�Tzg=���nҎ���x}/Ʀ����W��4�D��+��[�q��qUv���j��K��녆���ǉ�c�)K���E8��̦�A=�V�b����I��z[MOˣ6~~^�+Qze�̞��-H�aٝ�C��²�CU�h�"��<l��ᡞ�d
��"h�ƃx<�0A$�,r:�fu�#(1{tPz)^A+6����3��.%z�F�{�?�iPݛaj�z���q!�h%d�e)�DgDµ��g�LS?�)��^Y�/[}�4���q�Y͉~8�.Z��[������G�q��e8�Rڮ�T�$�5"7m�����h�'2~gR�J�$���������a������+���w�g7}T�APy�I>�����D���r</��X�����fn8xF��9b$'�WV&j3�<��~%������>^	��š�yI�N���ќ��iC�zL�m���0݁�-�}@�60$���2��GG���O/��i7!(�z��ĊAv�{5�]�J2����[U@�9���G?�B2��Z��,Й�cY>�3i���z�@��o �r��?Q�7[
�Ɋ�U�g��-�Y�i����2��,�QB\6غ��}l#oXA{�y䊷��fC�V"/>s�uA��?�s'gG��岁��V�%���Ԙ؋y�����v�~#@_�.�2!��_��weG[�	t>jeW~Q�:��Ѱ Z>L>rď�"	�7qڕ�k�l��b������e2�sϥ��Ֆ"�wx���C~;$,�i��M���X֌�̷��D6���A��g���"������vcϫn� �\!=�)����7�4غ�q���V��>��5�K,9�v��q�E1��V��b�s��;zo�-p<0v�=�!��M�e������0�v<W/���D�.�.�
�R}��nX�F�_}�Xp�}���u욄Ѫ��\�w1��M�1e��t1<�M�I�1л���>���W�\�����s�bV����R�|�������)5�}����TUq8�=}޴νE	��ӗ׷���F���12�Y�?�\>&��R���Ey�:_���l�H6_���;iF����� =�cM��K)����#6�v���*�K�_�O[4�y���,�e2�>���SS���l��w1T�JzA��ldmZ�,ߓ��>�F���wj���u���9���;��W�9�(=�a�dU�*ޠ�Ajі���nL���q��͉Hgr9X}cSv ��"�$��P��/�Z��2S�Ȳ9�	�����cꮙ�G��w�Ua2I�fF��>:�U���@��~^U�z�}Z}Z��\+��a�����e����З:9 ����h4'��ڠ����Y�㋈}Ɗ���S�� 9)!1l֮�:8�Ԍȓ�����Ny�Q�)L��6s�;����@�lK�΀��9T��i���XE^�xN��;!Q��xz<Q��L�.�q`�}�wz�)a%�Mz��
^�����-�n�0����������3�Ǳ�ꞽ�TS���z��nZ/a����f�?*�FO�]n(5���42���a���6s�KU}V_�=8���$����m]���5��� v"zUB��g��
�|�"}^��o���-b`���XWz����(�"d#[�W��z16t%�j�_4�5~1��Px]F��Pj{\��N�1�
�U�£.�T��Ɩ1B�H�V��l�.�d���_�4�Ze{�� ��Y� ��fG���M��o�4���_?W*d�wZjW�[&��,�l�(e�Z�h�7!]ew4s_�s?�ff���>�>����J�p�-U�R-��n�����j�EXA�:s�H�'U+�	}��ޥ�{��(@ڄ�4H��zE�>�L'Z#��o�+'��ܓm*��-/)�ܕ�j<��{ο ���Y�
�Z�@��4�;��#^�ٲ���A����I�&A+.^C|�S5�SI.߹���ۘo�����)OF��h-4حA�B`�O뻸p_H����M���/�gD:��� ='��{f� �w4ޢ�9����-Z7��v�{�tR�=f�<����Ix��� Nw�tZѪ�1��#�Y�n�&m+�H�FЩ��j*�s4tRg�`(�7*h��{�F�C^z���z`������H`�Ak��9[� D��^�F;�0\��`9=H��d}���|�_U�?�r}ݡ�/����y$Ke��uM�K�},�!��:b���>�-6v�;f���\��O��-
��*l���̼��~Ӂ]����G;�Nk��O�I���[haM��Mh�?1Ɵ��������%�b��˒�!\f��@�8��B����v���6�Q��֝X�Ƽ
/H�`37�S����F���5U@6JD�f�(Xj ��1)B\��m�6+]��l�!6k_��k8W�)��F���z7D|��G���eD��ݻ��*�āl�z�O�Iʮ��F��Zl���6j��=�^����8����j+2Ca�2n@6g��a]��!쁟igNb�\3?茤�}	��ir���;'����5�_D%��y�;�cF��Q"��U,
ǩR�.@gE�4�qw���x �z(����@J��([L`f���[�յ�{�k2���;.ԲY��C�������?42�*J��݊~8�2�a�2��'R�N�?��G��<&wb�����Y2,�$7EB"�@m�B�n��;}���:��2ҩ�ˋ�*�b�V:��M���8o�e$ɯO��	,.�yp�l���%# 8�+Z^��Ȭ'3���e�%�B}\��B�C��ũ�D|+��)_�۵��|&��P�O=�I؝q7Z��7g.f��$�)_�//g v�|�lБ����[n��ϋ�zC�'�**�#b�t�󅛦�ǢM�]%د��[���䆃u�ژ���f�47v���OAz��@�i-�"����*���c����V�ڐd�ѣ��:s�:�k�b2��]~����rN��Nz3B^����6ʼ�wD�����Y5� 3iX.bUۦ�c��,�ʜ��W�t��4��uS<�ǏuY`~��$y�G�N�RȤ��g�w��nڍ����+`�˚��fu��nF��V�t9��CXŖ�{��A2OڅL�
���ڢ/�D<ߤ.��lG� ���hy�@vh�]��yL��(" ���^eG⟫b�%�9q@��-&M���Ӑ��٣��@�7�$V���)tm��Aqq$�D�hJ���B���+
^�x12�P����H�k��Y#v�%�p�h�	�
a�R%g�����=B+����nE�Jr.󘖜�	Y���1�1!�|˒��C�H�h�~	����������>�t��()����苸���},~�
0zF ���eRc�r���=�a�!&��x($ˊ��y�Q�^:�
���, �M"6&�3����|l�J+���?������?4b�PԖKY�����H�c�3�XʴK��lUcp�;�q{�_^�gL���}J�Ft18�����;@��>������ {qH|/�( >U<�|��G�����D�KIx��sVh%=K�V<������w�]�O(S�pn7a����(G@�̧|��ϛI�d�]��7+!�!�qfv�*��{�����	�l��P �����:�-v$��Q��� ���������|BZwB�v���Id�VVEtfU����%���KE�ٵV]3�+8k08*{ɦ���ӎ�y�>".q�,�Q4��6+�F��O���.��m��9�Pa��Y���nQa��s�I��瀏THQW;RM�TYgm�I��N5�hl��'�n��Q>Cb0�hP����-6��/��ġ��eS�& �/��*/�^���wL��NF������-�'� �3RQ�R�<)�����Sӛ�kEY���Z֮q�����g����n�?��-p�!����x1]��w@%���K�vˆ��*8U�\|f�
{�P��h| �!�d��e�X��Y����E���1�8^���U����擝3Ef�L�u2�	�F�}�ֶ����=�!�-����"˄4*�X���S���h�@wT��/1l��C��35x[\�Ϸ��"��g��O�5��T�M�;����C!UA�x�V5m��k������k��ƴ�o���Lv� ʺ�m:��z-�j �a�e��<tuG�y�H ǎ`��� ��~� %�>1S�>�c��Z���( )� :gt!�i�k�K�m+�
2��\��ZY���t?��K4������<���
<��w��� >I�-**9�Z�b������~��ԍ���7dH�=���B��'��v�$S�?'h���/҅Z��+�2Q�����{i����x~/e�tp�e(~{{i�d9���Q�[��bz�+v�ۜl��Nt��2=�23L� �����ؐ�siS����,��kyo�?2��f\A�Y��+J�G�h>nH��*Z��uL�}�Oy>ܟ��;p��;�S���.[zS���Ț����]�)m���'pca��[��saqJ"V@��M���ܟ1 Y����vxz��:�z��Mv�T��
rױ#�4�L\�oϸ�<���:������@��xZKK~���Z�����r�<0C�c�J�4�B�Q�x��wH)� ��.�7��ن�ng�@�!�f,Ӊba/9]�x I��	V0�%ƹP�b\�-](W��0��^Q��~�*���(:�F��9�{��.L9�d�woP�TL�c*&�vx�)��I} \��6�y
�ԧ�I��R��`D�ݶ��� �	ժ��a	Չ� ��U�Azܸ�RJ]ʄK���f���8%F�{�✏#qJ��!�֔��U�˞��;H�Q��+_�E�8b!b&a#��""谚1t�w.m�
��PD�)��}�Y��J˕\j�4F��!�E+�XL�����aS��#�浂[*�Ȟ�!mnL�Y�Y{t)'�����n������	b�ŏBg �ՎV{��X���� N��jJ�p��H�x��'@1a��Y��ʑ��h������������GL�nߜ��º�h��&���� Z�3�R���fZ���b�Dl�Ebwf�K�JI�Ӫ�Fא�9�È)�>���R#�t�^Ԟg.H�c�<��#Y��C��E�bl���F���ɚ�N�ru��D���)�������p�r�ɵVȊ�p��N+|��o\I�������A��ͱ��}����ځ�5P���qn�1��x�����՟�0��W'�R�����!|2M�o-g��V����둅PR�WS�m�fO�V���hr�"�~�b�\�p�R�a���yi���Qw�)X�Xݪ㤱��/��u�}�N\��+_�M*�V�f�A,0)9��rHg�U�3.;A�!h�
Õ8JU�g"�9Щ�����2j�o���	��#�窂�28N�%O.FO͘,���[�n�Qc�z�+��5�Spx*Ex�������H�������jV��(����<ӏgO�����fjԍ�y�H�c�p@OA݀��3�p�#�.����B��}ϲ��B�U�4�<�Ws2q+2��o�Zw�gw���h�/=���X5yң �N�����~�(� o�/_����b���J�C劣]��&|�~^�;�G�	�;Eak
����#��}��xa&�4ea��$ u2�I�1	��S�_���7��@�م����WS�-5�OOm��������7ޔV�_P���r/�Ҍ�/���yĮ@b�^��~L�@7�H^%m��Q8	Q�2P��e:��\Dg+4�
�|r���M��G0��H��q,�6/�\��WWǮ>��Ѯkl,2��K�"��)�vE`B��0�7Z��5� �76�E�݊�NG��|����3�������B&.8��v�m4�;1;N��K�b=�� q3���y*�����K��h`�@���#=U��퀈��^'�)�"�W�,�Q�3�i ����e�����F��"����י�e�@�@����p�8C.�8����$���%q�r格��.��
��9��>z0n7Ȋ�(O�ƙ�N��$j����~	ؕ3!� �,m�&EG�<��_-�f�Ե�t7�H�Q�-�@9��V��Sخ)�Jv����[��k�t��![����z��Qi�ew��&���m/�T�b��`���O�hR��1��~Z$��F��w�~o�6Ɓ�kQ��HA���A�
�W;^���c����<�B<`d8�6<���-{���`��[�x��r���	�s���S��# �{���Nc���MV��e�b=]CK���.W��@�wIv��͟����PA�{ly���O�]��mO*v�i��KT'zR�Ǉyna��*L��,q��bi���Q�0(��-҉W.g�N���r�����p[#<�A)>�w�KU�y-��Yq���{S�S�&��1�%r#�c�����Li_VB�����]U�8_�D�}64����JW��!y=��� S��\���IK�<�����Ӌ�5��	�2�f��'���W���bg@��D���H�@1�@@^~�ۥ&p��] H�U��>�*��+��ґ�bP�:���f����J$0橕�93��(3�T��s7�kIgu]�S#PD���eߏ��g��+o<���L`V��@}|)]�T��{�w�+n�(U�ֈ%ܢp2�x�w�a"(R��KV�'%~��n�h�� R�L�!{z��o������D��S^+!��ʱ��@�j��� h��L#���.N��@�%�����4�ܛBDd6�~p�`�^����o���>���PĊ{����\BA�]�-�� N���|�4���
 ����	|��וF�����8q��E�~մ�����&&��?�� �v+����>��YoU��=���Rl��pY�IA���Q�6����0��s�d�������쓏�tk��#�b���B� ��Ǘ@.�kӶ=H�6��[uJ���L��8��oV�ON��k@|��>���k�����m!����%d�û���uD��7��i���>׿�����:���jR5o��ݯv4��΃<!�w͗���b�Ȃ��Uc[,`��B�m�y*�ߪ'.G>Y�8���ߋ�'4|�z�P	5>��A+O$]z�(���:�h�'h���g���`!i������e:��5���w�ɑ���m6�����&�a�4�{�cZ?�~&v石oM������0ʡ1b����&�a�<�+�����I_�DaU��F֗�?Ci,��l:ˠFR��*�?��qPW�ǳE�+Ǫ���K�
��	^k�1d���7�;;��qk�w�mc�p��<D}�� �_��Bt�F����7^��VY�`�f\>�2�k�<�)&Ӱe�x5K������LB��4��~I����պ���$҉���r�lEa��+%�J<�@�ҹ#H�k�}y��_^By#��:��3�L�g*l$���^m��6n�8(�����ܛU<��tr���h��(D'�J�1�=����kD�DD���i}�t��1pm~��xI��)�f�U�L���<��{�7��r�u"��A��D"�����:�y�Ġ�w�ΕY����Hb�?ԩ���`&D���no��he"'�'-�[Ͼ���<kYK�T��c�����)�0`�B �����^�F��.�y��#����c/F��Үj���e�|�}��	1��?+�YHe\�M��ŵ�÷H\X>9��%�f}�|�$����}�
��\t�F/�Z�K�����΍H�@ʶ�+'�nx|�U�dc�$q�LQ�M$��@����	�l/���nY���ض���ls�7b/r�Pl��X���qw����f�첐�W{ߣ�%�5�w/�5���ѡm`]Xxb 90��E>�D����M~U��#�-W��>�\��34eDO�u���$\�R��� ��9��m�q� B�f��ˁ�������sW�4_'+���5 �C��t����SrK~�6j�M�H�>$:q���I����2���W:�#o��#вӞP;bՖ�Zq؞�0��οV1�0�||4.!�h�U�����)lAރX$h�h��{YӐp)!���*�hW{Z'^�Jb:����߻,�=�؃��ȃlA�8DGv<�J��&�uxkVs4�<�~e�T�_����`#M��w
��~Q�ޚ��2\�,;ҏ��S¡��~\6���Ȭ�c�;�(a�f���$���.�A�%?�[v�5/�e�
����t����Gȗ_�@6=����"��N����/�������،�3���7.��]��F��g���H�h/C�w����$M��z�@�U����K,��7X�v����"��@��fN��O&u���
�Ɇf��5R�,�/P�Xx�Ti�>́O�hu�Д�.ys
u�=�#�ə��$y���0�奔J��?�̴�4�s1{z��^��xRS�^�l�c��O�<&S":a���f�V���
+�⪆���>z2 -���Q���15�c~�5�3)_�\;Y/�a;����t�)���P��Q�F�&k��x!ͳ���@^S�*w��$��J�|�(�s7���Å�4�����D�6I&�a=/Cw]�5�a���uV��Z�w]V}YF�gE>��";��f�#o�$z�*o��Ye�m�u�i�ls��\�?N�M���K���1ͷ�ߨL��!�+����j���%��%s>��.⑟�hH)"3׷��=Zz�3�*D��O���9�\�|��2o�vT��ƃI�$���9����"@���ew�lҮ@<�g�X2���6�����ߑ�o��Q�
�8���~�N�,�P�= �C���w�)�h6O�ȩ�F����!�0(������ӟԢ*zG�����Qt��n���d�Wi�G��Y��9۾ۍr/��4ק�|ǊGN_dd�`�ʵ{��8�E�g�o������J�_X���Q;/��2S�zݲzL��~�(�;�I���v�9H�Ub$��4��q��'�[1F~ۘ�`�G����/	X3�`jX��3#��|4���_�{|jh� Ǜ�1������"^Y�s`5Q�!-7���vA�� +gXOE򚅷"	�!gy!��K=Ai}��VǢ2߈lҮ�W7^����&'E>�ѵ���{��>�~��L-��D����J�g*��L���V3������4D�a��N���\XV�p
OF5��)N<���l%:w�'�q/M��!:$�'7߯�0��L_��׉��Y53���wR�3��f=�	qpP�f/���[����>�Q5?�*���Q�HR;h��>ǎƍ	A)1=�}F�$Nw,f�2�=&��v��N="��+qd&�U�Ծ�c0T7_6u�b#�i4S��!Ty�e�+ƺ�RNz4�׿P�|���5
�!�y�9/�m�_��|S+eE��OK�ǉ��/|��o V�t�`��B����w��SVw�4dh�i�NG��,�Yh͝ҏF����#��?P��V08{�'�qԧ��S�B7(�$�hȻ�]��V����o���
��]ն��k�Ɠ��?8��ݵ�+*����ݕ6�Ae~�cM�i$Wc���u4�GP�vN(���0��^b��7+��bM�mvD)�;�<��1�N������md�%jn*�ˋ.�1�ާ�]1!	��m�?���e 
��,��9C?�y��=�� �h�N�7=��T����nĹ���b����:a/�c+�uߤ�^BqT}z�
G�B������L��;h�,�x!-����t��!.b���oKv3�>gמY7va���:s��a#���6`<���iU�0�bS��+���Т*�A�~٬��+9C͚3,_�?������pq儡��ڏ��j�[	V ���d�	����~��|�@H#�u���m�]s*Df����fGj�xo2�+�ݭ'��r�XF�G���SAL��j�����}�O�z19s��h�aw��.D�X�b�=�4k�#7�#w�F}oC��IJ%�=9�pT]b���U7��ǝ��K�>� Z�����`mm�<����ԙC!zg�� �J�t�w��[K��ָ�B�ت��<��Χ���n�\#1.��爅�p�(C{D�	A�ʗ�%�aW�(���$�=�4��Ɩ��9ͥġ��3ـ� =r��������p�Γ闷��uW�6?P;����>�G���ג�
������J�kP�2�#�8�^#Gޚ��9��)��i�'�޼t_��g:Z��8�V��A@I���:�ty��@'N��1�.�zg�L�� _@^�AWV9��t�|A���`F=jY�0J�`�Jy��<��Ę
2{�p��{Y��0��`���3�B��8��f��!�U}�����~�A���g�q���$i�J�M��-h�� �����?�x�Ctm����j��{�X4g�ǔ����+}/���"%9B�uַ��&���O�;��7���ubU��q[�����UݛW�D���x���<��$�	o<⋬���'T���hh�a¾��fQ \4o
9-Y�}*�ܚd*���S-���f�
��VE����x M�8�;Sp���l`*��:sڷ����.Hv|����4Ɨ����vr����ψZk�m /h�|�XN��~�?�0O������4֞�h~����t
&�SDbն��%� ���L�З��]��fƵ	[����>R�n�k����Eʺ#o�G\�h8/�W�e�lU�(T�4�W�\:� ��`;>aݘ&��Nl������[ߡՀ��H2��Rc�٢��e�k��G�y�'g��j�0 �WIw$s�_�Q���ǋ��Ru��^���A4�O�+�Z��(�%�0(\�i�9?w��B!����-y�F;���Ŝ�^i�y�B5��g�0�|__w+r� cߴ�)�1��D��g̾"x�T��/[�Yk�� w���Yh�J�������HSf`;(��Q�
U���ɐn^� ��s�L�X�FD�p����$�e}���:R����$e��$|~h�����!�qn�y�h0/����<�e��Z�F� ��� U.���
�pMH"���߹n^߸�
����r�H-0�S�e:�ndE� !�
3���#ษBEW�4��6<]oAS�������
�f:��SQ���u���b$-�W�%��u�SC�,2'�{y�"�ݐ'�v)�Ǌ'D���s��2�[����4n�!.IWj8�nW�n���wss���
&C5]=9)Y~T����8=#8�X��0�1e�s�9H��q�bD!sx��'Į��3QT'���d(�V�y6���8���P%�:��௻2��R�|!�l�-���S�1��dj���=�P��㱧�V���(����m�o�UT�Ց��D'`O-WW����k����ÜuA�8�4q��ށ�)�fĦD��!tMFmֹ�f��v_�t%Sݾ�����"�(}��a\cs������m=��C�'�2�zc�4P�*�τl����9��x�"5�d�T�zb{�� ��I\$C+�mEn��2��9���e�}���ir�����g����[��5�*�an
��`DJfq��I�.2h�r�������.ӹ��@~��<�A���Ps�|������B����傄mS%�+{��d�h����m�RD�e�!��/��g���J�P)�8����p���.۹_!��a�B�3m��ā� 	���G!�h�nx��<%��U3����5(&r>�tQ���F�������J�d�z�rUn�c�4I�� ���ӧz�Zb$"�ԧ�$L<��S-��s�f�YM���<vǓ"���5r�^_��"�G�R�H<���
 wf""�>DK&��A�S̜�s�S����)�븶7�]�`��çI��,��{�k
~U�b�{L<������W��+�~�+׃���Ks
���N5��w�+���%����7�UB��#D��r:�3��;�|
����MR��SG�b�|s�^�g�/����7�1p����H�.�����!�hRN�c�V����c[��K7�S΁9_��(����_w݈BiYEu���C��B_�����;�ᑪ!v�|��>[�֧��L���8���1�Z|T��r}���Ѹ�r���p����Щ�F��{�"W�m̮E!�� �j�F��R�7F*{�����Q ��rӐ8�Mѥ�R29]�����3V�&��,����T�Q��Z�N#Ϟ�p���A��ԑ��IsԽ��Z�P�g�/V����9o
gx[LEc��ԡ
ix.*Lp��R\9Op�m&�%E�M:^ �����b�g�0P�n�e�B1���d�1Vڧ�"�S��-;�'�b#��L�N�On����A��`FP�'nA�bHا�`"��gk��[S'��&�� �#��(0�W������+$'Ea�(��k4E);��$�F\����yU>A��e�6�[�؄�ї���Kz�?�c�P_Eo���u�y�'��#����N���S��p���(b�&2���o�A��ǽ0+�`���N�?۳\��p��M���J�.=�'K6���z��CF�@�6��_��e�?��y�������7�(�+ �d� �_Rڕ1�oRD�����8<R�XQ�@��jԅ�m��lwXYV��U����'�ȇB����\F	e.�xN�z?��6	(�J� ��-F��r_S��Ѽ*o�ׂ����m>CV�/%�l���§������x��L6A�Q����6����wR��\���2K� Bjj��oj�u鸚+���g)tND]|���F,������)��#X�o@j�2����?�I����]wH/��V^_(}���$^���V<0ץ[�G: z��,K򈶼�z`�|�'/]�kW�/;tӜ���jTt��<�����b�Wm��v��ְw���y�����2��������~��G��\8���L�Cd{��5��Ɲ�-V^��nzs CR��'�Qs��
���A-�������or �p�4'�D�Á��N�lX�� ����#{ �s�����3����C�i5J�~i��\G/��@�����(��@��l��;×���c3o�"�;�r����t]�����ɂS}:��پu_��c$�>��H�d[;���S�GS�&�q])B]�|�t[m�N~�,�!)�dTN8f�S����ܲ��5Gg?Fk,{Vg P,>�ҞK���Vy��fK�[0�X���7\P�BLN%!��Z[8e08!3��H.����n��.��Cw⩍އ'3آ�4 5~$&�.� ���>u������kcY�%� ���>އ4���W,K<j�Z�o�������������S�� -p��=��)w�f੗����>^�c��ܣ�W�� e���l+�֢�u��R��$!U!��ͥ5|=���(�Gz����K�"����%영��6���E	�$���f��.#3������+w0l@}[��N�E��&f->1�����6���GXl*�zI�s�`��u+���|�[��LLT�0("��k�~E�@������wk�S	BU:7�5��� ��>i�����8�AC����Z<����6�K痛L~�D0��Nx��DU�G���ɦݓo� +f�R��C�"��>�����]td��cI��?B� Y�L*l�\:��0(Us�K���"��P�gVz�6��M^�;}O9Rǆ������>@�r�Y��=�GC���_�����^<���x��!n
iVJ%�Rd�������`[�_��2&wNY��Z8X1�Q����uU\鸨#J��Ze��Ϧ���_�窴.�l,_��t[�(b�kS*��,�b��/��E���5�i�����'�R@E��QO��Dc1#9+bDʉ�Ric�L���d��d��e+�td̫�Wt)仃�����5�^U��T���K�~w>�͓=�5^8B��ֺ��s�����c>���ၟ��MRQ-�n�퇠�r�|�hk��	��Xx�3C�����o�5%���[:p���#��rf�5�a?3b»�K����F��E�.�N�_�#�T4� ���3ʩR��r�i!�UX��$�u�C`���卋��\ep!����׆��z���D�l�C�^�����D���>ʫ��@G�ɨ�4f��X�����,E��:�,���˾����
�A�}q�2��Cp��Ξ��XXKZ�>��\"1��q�g����PJ���-�@IF�Ɏ���	
�M��07�8�	h?���sE�>L[�9:8dY�ke�W/���	sb[ƚ�M+y���@Tf��O�%]�)�Wl�8�qF>P�[B� A>�7�.��9'�u�B,����I����e�1h\��b&�e,���6!��ƒ<�������`�<���\�O�竓X3��_y~��ʹ26�3���g�=+��啂♩�5t�ǱM�$Һ�4z|~�4q������s��0a	л���F�3V���v���:���Q@<8��w/�F%��U;s1��cu���8��WK�����]i�o� �b�E���1��A��3+�cʏ�بY����z���ٝmv4(#���)�k���@3�/!���6�_�
��M�G�?��6Ÿ_-��~����}�l��ʆ,��u��9w&���p���q�����@=�9�0�3Ȼ�����i�EZ:Ş�U�|��)6ȍ�5g�V�|�,I����v����@�u�ȩjf� {�0>h�h�n\�24�n�;�3"��Lm�>��&0��/&P�O�Q�׀����w�-�|=0��2zŝ�d�Z,�w�sb;r��5�qo\'CJ�~��ͥ-!��^'��v(�����-�	��1ߞ0Ӑ駵�%wEpN³��}����Ztk^K|�:G���5��qc4y��Sd(�Ǻ;��m������!lM"R-vs?�n ��,����t�w$�e&�����>ǯ��{^��^o���)5Ԁ������*`�����'=s�t\�7��l(�21� �e��F�$�L�	�7���ˍq���v�X�C^�c2�^� ��\��|P��J�L�'-��2�:�B�����d���X[�\O`8�ޭ�$�Q��	U֛�PTNYF'1��!��zѰf��(1�ZX������KD:�B�2�(�H��bId�qj4	k<�8����n��`;��K$FlV���)[z�
�?KK5�~Ϊ��u�|/}3���VPl+������z,D,x�X<H��xժ#�`� �j��5Jv��l���=>P���N��dXdQE7��:�'�٠uO�o���E�NR�+P�*�L�?K
^�)����}�m�<O4e���Bk��є�"�hx��X�k���"�U܊֯R[	�%a���Hs)&��)PC<�:k.e;��$�b�5��$U�qō�o1�Ѝ��{&�tU-y��2�V��1�p���+��=~��7\&R���Բ������]�96r0�J�#��t��d^ŭ�]*84�n(<��9}+$�x�A�¤L�;Γ�hǹ�e��|:�3�^��%�Y�P�Dه�}dɂ���{^k���؍2����ɟ{X�H�*�׏+���MR��<���xeo�,��Κ_�!��2�Qۊb���P�m ���ͦ��&�P#�xڷ1c������_F�]w�/ۓ	|�.HG�jj;���ݲ��%�=fb�`�y��2A�(�-����o�!A�$?.�F0��da�%&�z��,h�薊m���Y�{h/���\�Au��QG����99'�Z0^��1k4"����ƙ��@�IŸ�1B��G�����2SS���U{~�^��6�m��'��\ӥN�`˨瞱x)ۂ�N�Z�����J�;�� z"�~��*%a`���xَ���:�� ���������.%Zȉ��;�
@H-��T�e�$��^s�B�u���d������q1�H`f,�\��
�� x�V �ĺ�#�,�"�K��e��LUh��D|�#K��78 ��0x%���4������,�Z������FF�H%A�L`�"�c��S���(`�Cj��	tyɘ4��*!d�:�<��"�\O����{��`g�]��O����q4��Q�KJQ�$�Uf����E��peo��.��������������Ì���lZ���^}�Z�� �,�J.Y�T�F ���	Z�s���$sC���fP�m�-�$�Ɯ���v��t3ה��5̏y�_�5ؼn��ؒ"`��v�<����֠6�բ��/?[�m<��[�����c�^P� ���G3�=傻`��}����~��Pں��g��{�I�T���E�;D7ul��� ��j��7��.��H�uU�9��ќ5"X`�������|Y��2�^>@+\so���o]�;�=�v���'.�m��?�Y
ƺ|%����Ws1��%HGP>l�j����/q�|��0��7�M@��M{gU�є��o�d��_9��&�Ǜ��Ɏ!�C+��u�l���S�7k �ɜ
>��3��W����;5$B��Cp�y���R����q
���2[�5ѝ�m|K;Ļ��$�D}��ގr����uJ�"@8eܵ[@�r`잚��c��� !�����L���_����^m�KF�zC'�[#DU���,<2a�m���{����M�{�9��i���T����Oat+������Q�m�ɡt�hI����Z82�1�n���L.�O�xs$�NK�<��rH���zyx��m���=/��xK �w��K�����%zɦJ��yT]xb���w�G����I�L����m���D�����r;
w�N#���9 9����i�y������_2�P����Ր��y]�l8�- g��]��1�(��~6��/˩�8	z�ײ�F�E�F�Cc73��8�x�ť�E3�ֻ� ����(h�s���`��ni�ʊ�;��y�[4 Ń��wo�s�_|���Yݛ߅9��j$�-݀��ň$*�n	W$vO\���씕S�d�愈+��Y���Z[�����:b��P@�-dx�8��آc?K��m���\��"���T�e��ac�F
��B��9�G�x����z�w�a�ߺ�Z�.H�-�����i�K�������
=��鈅�C(����^5�V*�Q�C;~ rd�n�j�_;4����G|�D�ʃ÷�`t2vl��f�,9RM})Ҹ(i�kv�|j���G��/�D�aq�wN�X�Eȳ�D�͎�����i�<�1�m����LO��"$>��YvŘ����ݢ|3�>�;o k���4�{�|s)X�Ǵ���c-_�m���2m����-XY�b�C�tJ�po��NQbIA힚�Stj�KS�W��Ĩ�r�f6�x,N�~�%z��{��9�|�$��Jts�Zd�千<��0�������."�X��"g��L�_���g�Ĳx�y&��2[%(�<���w�!�W�}��C����礞3�eQ����?2�­�x�*�d�y^0F���] 0�Y���2���u�-}�)W�#�y;�d&M�g��j���g�����\x���j>|('Pnc霮�f[�����/����/��v;<���$�Hc���Z?|�F����m�f�a!�h[g��U�?Q��