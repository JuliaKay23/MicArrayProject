// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Hbzsr0h0OtjHJNaLuy4OOuXeakv27BDJ4TtGXsbi8+9CDpCZ1wuCaNjLpytCn4M1IwnGMtuwY1p9
uMQ0inTWXlnZ8EqAqwNVa5Ug0uOVCtjTLYgpXYwtSrbQ6SpAvvRvJSpZbSdyMuKqPkXlbdJ3sEpR
wqJ59FFbKeX/MBlmDghEJcIYORi6UokznZZwXdXr5nHfJLgYikfVKpHY9YI8R3I5hIQ542Mz4Eke
KtpaBqiG+KaXbi1FVbeqD0EG7oabEx8+9sAdDTQfxywjT/aV5kWnmsEOUG4o/o1Qs+h70ZinUmV0
YWBybVRH28TWCecxQ8DCl8VjgDxZZWOW9geylA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14000)
myC75mPd7Om//Y7PbvQsR7gGEbcoldset9ZpWfmzqmiZj1TuuaR1mTpilZUrBNCzW5wWDOlWXav8
0YxuNNrPk9pA0TKsiHQjpZzMZUhmN3n9RfhyIJlemdqbmExyUslMQyQLzQD7lwj3IbXzuH7k7LPd
PZNDvaNUeM0tDx0vtD3K2bqg8p5L8DsmggbKjZHLAExJuu3p9jZrXxaQxHJVBG31Bh5S7eErgAs/
KGJWLKevkje9yE+JkH0eKYev7jQT48lOyZ6B0WKfW6eVuxfcRUsCWMTfhWKcMKYPoUoIVAutH/j+
FSjp20srYmaUIlGbegTIsPhDmtvkhHoLaGXeS4TK5aXE6BJU2fG8B44XllRglbF5zHgPEKacY7VO
TxKgAimW2Cbj0TDE45vhvmN8somblWgb/ZLmE9cRLbqcHbKKqAfF3GHMP2PDRBL6gsdbq9K1EoTg
Eyq8CZ1/VSL99ZO40ZRQ13F+O+g3aui+Xa19vWwHAZd9UdimTXtdI8Rnsxc2u0MK1k+TkQuU/p+y
eRwGz2tBM3zZo9xBp5aR4xzY/naV8btmooWDTx1prkCPKatpBtRFKLpXpzwseijkHxFbS8p/qLyh
zMcPcOJxIX0vJPhDoTTR1oSzmNh4wdktsXGM2spWYbUtjl1yrJjPpdj0Fl7O0mmoMSuacZns4KTj
Kf14bMCy5NjZ3f2Ok2OSWh/Gl2Zizp+S9lll1ZeUJVfbZ0DUwDzSLeEWC9FNWH4990fCVdUBXHDB
62JeE6mFY+xD4nmg7c7Xv7v3iewm6yoVnf0kAa0kPhMWAggVl9Q4hN3lK0RVfUhAyWFvyJ8h4c2V
GMWnu5LNcrHF7AfdR9QzQUGjlHQazy4KUEm+Om8wxH6OnrotAddGRIcNIj1quAncD0AAMavxxT1p
P44XYew44xUnHpJUmkts6gOs6Dmn4YIkHpJSn0325wmhAHqIDOwLdizzRh5cEj8Ilpd8xj7/hQSW
OeOqiLe7nFAiNDb2O8RZwaSd0r2zDayhgYaaUf9Qhpm5RLOecdP+zQ6khxA2DSWqAirN02bqvI1M
Uctr+d7bvcw6YLZS5MRiU5TS9ofQzzrVAe5nLb2CM2NJqCthe4m+YrGSkJ1q9TyfCBqoKdIj4FDR
GuQulD43G1ewTIpmUwhhc0RkvBYT06+STQlfbjqD89p5tFsdIKHMNWrBthV1S+HJuWr3FzbsI8If
sh/m+9+aC+fMjdv9zG+A5Y+tDshs9IXkwmX8qFaQNcMPatql/bLBoMNwJ18+hCV05t01SqYyadzQ
Wux+T/3VXntsqgCGzvqMsQEL9idFwegMn0V4Ruh+fw1WYnAeToct0fJTjQFHAnfc6zrLKfulwPTe
3MuUfjVjPUAZG7RrxDwJwCw/77KO7us5hmn7jPunQrstyuecoVtc3vTeslC6lDu1bCEMt7tFDTnN
Q4arTz/ucym/I/jYZ6kQyxxc5qJ4LFdWvEhb8cd5/cwb1wpWTLE5XP+wjiiZMTMRuW17m42T0gyQ
cmVX4PyfRTA+oaj/YPYxzKPKmnvlJ5DEi9xjidWA6wxGXwDBmlHluXUYNJzzdMngyPhX57jXwl/1
6BLkpXXrBTPcVke6OIwAD+ddTZo5pFp/hp3sWQtbmEzRSgrzrLN1q8WxUcjxkAnAkBvFamJ4hZ2O
ROqZXOEy8ujXtN3bEwy5fKe72e2vnwpTD1JXg0HOZ86bS66JUqx/FrCDK+oNSymqhmnG2KNo6cP/
fTwBB8R0q0gV5kUdDTXWCrC9HYsnd9bq1cLBm9yRpVNRwP5WlnnNwR0PUxY8tMkHRwTuj1VsrL2r
4M82l80F3Hcf6fWJMQ7R4F97i/8oKw67WtPj5gmbJkx6r5aHH5v2ZRtp5ze3VcDLnFjSj2DAHMjT
iAwWCzvwHBA7VctgkzrILKO4PjRARpM/saWXO/J0stXpC8rVn7tAUcFdrBJLg2VwvxjKM/4g4Ait
fE7sMKbDwJy31odvi6MrNg3V09BCWw7vSCvoMqvgIHuTb5iIqPJhxQIkt5heUzRa3Tnt07gWkUjJ
CLQAUQEsvCT1KiDDFdFR+g/pRJr/sC3bztgE3hMcuVwUCdqmbFxVL7bpYJyIlVs6IBKKZSrOb1bN
/SJVSb7Vw8Ji6jm+VMi61N1x4e0AMKHTCaXE3DrvBK5rqgXl0mTz0TfYNTZ+k6gZt2B7/hotAZ6q
thzfXfcVrEblGMCl1j0LPxswD2WomDfmjb5BAq5bIXpFyelSu3O0FlHDw6k4+IvdofW8eDk7h9VN
+G5GL3fQpNFYu3ELaX7vbZWctFhaJaMsNd/a87zUES3VnrakYrWCbZHDfzfMm0yssQ8wNvZtppwt
Ps8mk/EUTp4nWzx1yRsv6KttauK7nttHCcftIYiFeNHdyovCEHfgCW8MhQ2CVU3F8rRve6oB3hu2
GErDAM4SS3+ToU2k/YkqxvpsUf9mHPmw8KtFXTmfbvNCT4pQe3tgAT4H0i16mkBRDs40CYimERP9
Q7aOlCOfH9RTnMzGMy5rs/F954Y2BJFHJvuzsrHLfrXn2xMznZGz3AGPvec4AfctONt2Si+4VT5D
tg0WAYXhwCSXUzCCW7BtkZlAwHlx/61V5KjwTV4jw0TRb+88qQ3fA4ultQtdwUgQYdRQH7IdXdeS
v8ECk0lp8RDW6OOxzq2L6lER5g/L5sd4GJC+CHbRt663RY6BLtzcqxbF790hcCqDaO6Bb1an0bJ4
dMw4+RmE+4q8Mb9Yw3Qn4QAxXAlB3pnLTLU9GUAdapAF4JzLPrIqbFlF8OqMQV/NLNfLsPlLR7HY
LqF68DNotishnbM4fc2W8KWTAzOeXK6G3iEmwU8U3Esdap7tMkJOD7v0xTiuS0hAI8obAgWR757s
J4ofwpD+23KNg5T3L3VOAnQ8mtNueRYvETRqVi7uzHwvvaSzsFi5z+BNXtOiOTOwPNdQwOkDWjhb
MjWJ55fKQypENN1W7a2qbiGzrFNRAZ7Vu/Rdk2OY6iLbuOkh2f0Adwfry0RcU7pg3Vwlyf27kl/F
0Hf7o0jQoCcfB+8sOlSeHjZKm/jskFiaA4NjV0IF+QzIcSFk9RARmpHt5T3HGTie9vrcUsaXmtH8
yK1pbSAbXx89ELVXjGYHaD76nvpgbsHRHMgSw/lYTnOKAAu8N3fIg6UCfh5VRPzIIKdABjYlfnbC
E6I40C8Q/HLcvMjclZ5kx0b/ndlMe5hjmnD5Le2dfFEjtio/NyzY5FpORKXzQdm9la1lQ2IAxvUv
XmBs5gRxdSqOM+V9dE8+B+Km3MDvgCHJVZ6+95Ks1N3G7Ux5CtGkOxf82RddsWa1OkZh00X2yLcC
0Mwp6+EUC6STB8WBXPp19d7OjdeRe6LwgR8mJKMiVSZ6OuVzmKxtW3n2OFbXm5vwsDJH3ZU5Ri2P
rVfdr55iWp+zdDRNHLdj7/neXxKMQK6xvPQ21WcDf9V2mlz8CluBuQYVQSrG8aco3go9TnzEsa3n
XJ92jei5xy5mUkVygn0AiY4J89b8nRC+BMF4Il/PsQOp3Hlk69S1Dth5M7bqV6YqCFilYFgI6Sgn
kTSiN8saWAAo2JoJflp/xTgKsmzSbECv4K4CZGA1DCqBtxtxEeCKCQ6vLo2rJ8ZJ49PDZ/K5pG/s
NgWCSWN6ez42W60vUCoYAcIpq4Y1H8qf8W3Q1SUaVa0Sw1MWw8kSmR/7hqti8HukIwgq1XaJp5eO
RcFPjAnFWrPD21nTWwRQnyqq0DayV0V3GIUzK+CutxtD2f4d3TKxvi/XXQrWnlNj7RY6lWDvmq1L
4qkMKpeJoja0J0gnjU/17LTNMbVwkBVqL+7tfUhMH1y8FdmMoh1jBEdP2x0GVCw/geyk8h2ufh0y
lNUHRqj+VxJ++46+d/w1VJyBTVxj6mJhiCpY8V8nHI+jzDpxYDdj3afVykCT5PjjqLv5qbiPIbOZ
HxXZ6eP83JewQxc37zp4u8D3ijLDM5aDaGixXQWls/qSIf3cZz9PgLkLJ6GgeidXR/5D78DRE42y
2cWOzT8KAFI1GBFeZ3vj6Cmk7gyhjFLIsQLTWoUFxnBUNA43ZCmjqXMsyTnzaoPRzcXaseEQTuKe
yT2ySRWoY+UqHMvTZdBGYclULqwsavD21AYRNewDO0fWkxGH5MrIGjNYi+o6oRtC7HDe9y6YW2Z3
Rxt+PtI7U0V0A6xbshHPmKJhO/PPBvL16WWAJHETxqcBfgzC+W4aNYeByEjSMzuk1PloOlf8RGEm
D+59+appjV9ByA2H1i99RXFoLjgZMUrjQozDDJowDyZNrMQkir8i1zuJ+c+VUIAt6/faZfXBD51V
dwUxZi+wi9OufargcfCtKwatgArhAJ8WGaCcz8B/L3avVRQMJLo5qB4w1StfM4ZFooKETTsEM+b0
dq1VoHAbFKsrGYi8ZsXOROWI469Eu2NbEPRxiczUHW/hmRyCfINbZj3/k4JVPVKOjRa0GpLqZHtx
yjJzq2bFQpMcfxnF0NvczyVkIAi8yEcQqctgb9o9CbZSjxaThTQX4twKy6cBsu0ZkE58VZdUa0E1
nqo9dmh/JsuGDbdolrUHtqmu3qDuAOf9vxYOdneNrsd1gTo5oujI2gdOOycOAwdCAT2EJTwBHWM6
Ued/F69djrgJeV3Jk5M0WXSXal/lth/cCD/djRqWndsBEhtmxPEsd4cGlnxFK/b85B1N9d/NJ++X
SES3vvilCzJ9Xq4ieL+kj9A2o/lLOwvaGAXWsIjsNA34Oa0NAdxWkCrv4v6GrKy1kpcJ5cXV+Vnb
AZRtc0yH+UKUcsA96dOojFBs5tESkOnEHUJ84qBO4g5WBu+oelmTzsoMPmjZHlcFzM9X1+lH0UXO
jnWUa2Ioad9ntrfIk63gD3VwqWbpXJQcqJ590PrdtCC5UxLwJ6cewz1f9n5HOmGPDn5nvZvcRSfs
hb/VoqNnCqU2jfdDWklF36LtZkwlyqDiGra8MGxYa4EEntnhNFUtIo/2pm0JsfkFD/augHjlY6qF
XWIw/wO1va35bTh7VxbJ8E2bwUbQrz1hPP2ho2d2ZYUbnS8cdjPWMj0kNYcrt5jeECRzA6M5xI/q
sLZVqNZVhsLGYvCqRGFCI9Y234wRPv2WutP0/JspZqYMovSPNB2o1EQN0jgNb4a2QhLV5VLywf5l
9i90JWBaZpo+0vfH3s8KR11jwQpY7/nMxbE9TVQucP3q8mY2jhW/OH4moo8yHkT7eR5i97+yByN9
7ymWazoygaCViyepekWUMjAkiIazhy0Nudxtl2T2Mob6n2wDf4BSnc4OfXwiclvtLTqYt2b0MHVd
xJKZ6mGzldSIrcLOrPBPmhyjMmCRsIMceW3SzwBXnCPFT7PzMToRGG5fBkzSOyWdKM+a3Xoj9pEF
ayAn7vxFATcMckthrFn86VuYaEo8+v6z2ASnUoY+iaNT2TSwf9IpcDBrsvDUj196yIsl8SEC3PL6
YleWNgCwgovvS5XNZP+4onbBluVNbL7D08wS15dRprn/T2ljUq3NB9ndiZb6d/iGss41ieXjLl8M
QeRpCeSzPRj2ynELyfhod5K2924mhlE82kMT1vyWQpBbbAvDflEPKCPfEM02N0QUFRXKd1uHhqSQ
/9DdB5TL8ZQFXyfmY2XkuwIjyD7wmmsjXqPcMk2lSEoXfV92N6+fAFjJ5VvoyQvkVbwkNGWxyQvC
BMkBZN9hOVbfdulVXTw/n70rQBZfbN/uB6Jd+nCwUqTEgtyXJn9v4iRh/aCD2maxC5EhXpkGMhSa
4zh8EzJsG+xoAw6la6G8JMTudgqFBODfvrpQvKAnNHZrrR0HDoQtjfc9Gp1zmiOmN75vkJA/94HE
1NP8Bn/AHobZRZdE7RN7iM2pmGnKFoSjeiZBxErPrI7MpYm/MQh0lCthybPCu2vBwa8TId71oT5d
sm6x836cZMuklrcvk8Rfb44BOcaaX3MgEPUYV1S9g6+Dp5aSYISi7Uqy2+Z71lmTcCdO7uQrifJd
HDzlXdA0qhP1ozADimN4dvaLNdNOIH2U+aKMqnrUZTjnnAayM9D3H25+ugz81DxNVJ6zliFVI+nv
eo2mu0AmbqLHXbSkCStAMf+K39aBgm0Cqmhg5vWehM3xRExPtuaTpJ0SYkb/K+4zmmQwK62MNkPp
uIdVNe+YNAvZ3HmoM8KLO0xPlExPMsgVMVbfTMETCk5s07YL0GQsridf0EdUqR10yp+ktxXlZOMO
NNLo0JGvgERZ8/oc+MrjNWbJPh8/HVAE2bR8zM6femKGUwrtg5Q5I30L7HRjyOO//rdiLupaLwd7
OS48fqINt6ajcspLXwfA6ku+zt8Conz2pgD9p4xZttdS2j8A+6fzBwn58m4YP6noeiQJ3RC/EVXi
RL9pCrNvFR2/kPuQ9taW+8ag94ZXcAiA2DrYG57vjBXExrblkQuS6jIFW2O0+UPzt1nAHX0MikT1
YWW2PqxGa6FM1U2BY+/HFO1gzp0+6eLEmdi2vh2kbg1mUs531MF7e+puy4yD6OUGDGMDYK2HSGlO
2oHMqH/EhSfPOicqbKr5dqeQALUPhEwRS068U6IvRYARDrjDHYPZ+cdVKgsxbrvEGyS/5LoVj7zF
qfI2P7GMqj/0oH6HQg004XzdNv7h0Z1Ka68zpuZoPc5t4xrCe5a54WWsXlbkjZhtf9Wn7vmf5Fm/
f/Iy0TXcB6KPVa86vX7iDo1FmlXPNIGNhIrq1dDwuVZsj7jS2xfyNJS1wk/UyOU/GwBKwRPyS/aK
eVPHguwwUYdkfdMf4fFVP+D2fhDnAgFlp/lHUU8h/iRt+ajq0a3ImUg2MTnH3OzHecPwxHrzG4qv
8gbTqNQPRhpvjV8To+Ku8hFjOOd89eTMUAKb7tMLzOYsuZYBhwAWBH9wHQR4wCuTtaNiVMJLDAqK
aMpaBuYdNcf0DlTPOK+MET2apvmVM+yd/B64EMGkCNOT7U8x2jfmje9NUl3rzwI8EHHaYxSeGG1u
RV89eNTGO+9+oKmNeHFNZTFBL/T1e0NUCcSDzO3zVPXCETO550JfCfBkm4k4jY3sLq46w26/4+TF
mydeQQR7hbAjWc6B4XsxJIhDRPDREnEn8gbsa2DguFv1OBXMyTIWq/7/84aySNmWMe5ktQfLjY1y
so3wV2yWU042S0XCMY5TaEQV4tdgtINeogwinfQdxCq48UBaqG938CYHM4Bc81lSsfmoLcBi1UTE
QW0tbjNqMvMeg7KliwU+4hOr+V8ejtxYABCDhu2AbkjEoBpPSYSDVzzVfErzweZgNP0bxft+Km3t
88m6ij9X5LogkE/fq6RZegkZV0POZSHiCVTNxGHKmedeoIFHlH+UjJ1kPc92jwK3mo27a1U6CSXz
kpSXyNXrqHnt+qM72IsDlC7YmXUqWceGHFwVToLotzKqm4WKPp/bF0REmkCmXmLRpK5aPAm+sHDR
PFJ5NcGP3PPHWiqrnUHxEH2xkEiKMQNZ5rEmSh8lOYiGMSzJ/w5Igg05lJ0VbcaQE5kj60i+De3l
P5V6VMcWvn7CANeck1/zDgBQtnaIzGLycVKfvf83KY20pdEq+snvl31zIfHBv82MGrwSqh4ltVat
aPv74oGv1G6yKxQ/ExE8AIVf4ip/WhRV/G3neret+OIZYd+wCK+Hpi4NC8z+LzrWfGo2pzxCE1ln
jkog55+jN10sTyG1LdhrwYeyBmFnepO1ceZrHjM4Tot++/SdMo1Wnd9h5CqPxrlj1mYvsamFdn+z
6GU4fQ9JC3CsDwhV0kbcKDY0Fl1IfVmrZCF0LcOu1jF23FbqAEl4PVgddqfMbB+MD/BOGMmdLdIP
7rl6/BbF7g8fh7Tq2eJbKylvanUUow0XOIiLK5LyBdCMc05DecJu/JYfVwHu9NaXaghG+o5oYjtP
mPgzdLjmeA9nByked0LDH43Gk23OS14z2zWkbjIS6/rhVq9Ixpthx8UCd76I2NneBVjSK8BXbKQ+
VlNlq8TvLjmmCap3vWEpkjodeAUQvBRc84qoWynJnCsNuQNR7U9BnAURJFKF4L2cT+RLR6+ZTwyv
sgxfncTUZBYk+TaDzRFDhYa16cL1kZCXDIPmAt15dtzmp9MaaqDjL3iUc2LHVj441A7BPE69fiIw
YSBVszehiiyMs5FnQOvVIAVA9d57m/ak+QVXbGNl9ZigG+DZZB3pAKo+854eeOIKiGCpCMEo4RUg
DZ117onKahWzEXXgoRb0PQFlyZoEJo6gfkpTqt0rywV7Y0/LNIPKJDwJffevWKdewzOYCFANQWg3
lzWpEVXuSlD+UD5S5Zzu1j4VYmm+VxnZ3l+0Z90+fwc+iDfvTzcMrZIfgZ9ZQuq0wmY1z/Z3AYRc
Qcjnl9CHzNbcmqmhthDoj4FOswaV6LRo+kb8MaHkFl1kINBzFSaNOoYsjwMTL6i/bid81rZO1mXZ
nlgXtTepShj2t3TmntEE0wUpiC03ch7XcVHfdYraQWoQZNirEAMNG7le9ioRP46+Lh6PUF9J7Kts
qEiEMJFaodlht7Xo976srkcT+0cvG0hFfsO96yw48JeMdzmABY2SuZ2E8YpsTCZuoPK06ytqXFHA
+M6o36mFi+7aA19iMeg7n9QlTGgpoB2dmnbrowbGHqgoOFZpQFFrX8+341x3vkr6XxQlvPwIJPDd
nOnPcRbUP+sxT6HGlcI4RyVZfDYJUd7JDqNlodH0iXzjEJyakR1vRzmIXpRaQWS1DsFAjV8DAE6L
mXLKjvkdl3pUFkCnDiEaWbP8ga/gHELip3x+7OTYZWUidDF++5DjItiLDDBwIS9krgx1LsyC4jjm
MqUbJYVQlaup+C7iUGrY8VLAM4kEwyzLlre9KCLGqQ6mwS/2xLrOR8ggLxwf8lfRMIx3gS0mgarF
Kl08G1z1rgVNPjTfF/xbABRZ+DL8q00OBvP/RH5taKMphsJ1TeAHrNkfODI4XejFwkhdIq7+lv6N
qQC/GwYDJnNVhIwdwsFrn2yHiNGSjZDJAuokz8keO2taStpsbhCIrBUAIgbQXXzNxF0+4nm+cOpM
CmOeEL9y3DGF7yDX9AZrQwgaDfHnGZyP4DB+M6TuLXzuBGGPNMHi0iy+z9/ZWiY50U/frH9UlX8a
2cuJp1bIzKKMDVph/2ZYdyIJUsm92hRuDH2Zl/kNJhpNvfPQ9DCaGmHqRDJkUCQDfKpzqI0neP9q
9Tjc6t0d2Na2k3q3u6aj2XnraeVauzTmK+7Bx7wZ/a0pD4K4rCuaWbJZwgwm/Mkr9e192UBzaeuf
SQgzXmmIRgZt0DtCiQzjvgb72LboaCDlwtVVR9JsGr8Ht+vO8FgZiiJQHyn9Whjj2QnvfwgfN9tF
qLptE6i+PqRYIMit8ierkSTabuaMupPb0yyOqVvVBzXf7gIQlhJ+Q2TtOodAV8zlEag937AkFaDg
xDJFH3mhRBe7CORAMZFOYK6C5lPlDaVNpRmcQUvOd0R/5zAetLlwPfeYbqNyTbXBl781qLzpUSVK
UdzV/Uq4DUjMJIRR/5dAcwxsL5VJTVSi6M9OM+wfWXSbw2PXXe9KasAyBI40RNpSsjGXPsbDmd+4
8GmZCpPRYblKz3QAr53smVUfOfRWBHUKATpudUSp3PEUjSsvH5m+4mnbDGT2bZXAEgr1iGPpiDpa
Zy66Vj+efpv1ywC+p6IJGOPinP3CeVCwc+vlcW0KXzhASDm6jv5tNUF+6L93+Dgzo/lYd8VsilVn
eIGfk/0bxUBncZV73V+PnBm8wLYWBRxr1f65acS+xW5TirDR8jPAhdlhZAEdYeZ9Zoqg1C1/2/2U
tN4XLWFrsS+DUrRzJeJsfeeUO2T6g//G258JkMq8kWrC/lUNEY8xqDgt7ThusF+FX3WvJSVAT0aM
QoWWRbKFH2rwaxrtqWAZ9xgZAFPjMhZrOLiAcJpThStODef5AlfpzLnZPCs49wI49eRDQTYbJbTE
PqJ9h1UCoGp/EmzXR7wk32IqFiNOs/2WhU3jDbAKo9IlVpYwDVbk8ygJXCpbpFa4OLjHfAI5fw21
iszUHLEVwdhEyVn851WCcXZgnYKMwY1xpSYsNfeU7eMXYm4i/vceugkBQSkY+3cNajuVs1wfCvPB
YnmMX8R3YUdKILU5x7ZWHSnNjQUgUmK41T7Fjj+FRulFXzuv4MYByVm9J/MsU2Dod/5M0AqgdrX7
w8nflwV8eLjGHxySF0YcKmbUDa41F7BGENae7gQAjHEtv7rShDMRdlh3w3M/gJrrL2tG53/3vGsl
Nvz0+q0eyZ2XHmxfFw6uEMfy4zeb4VVRMrE+0B87wTgcDlQuSwh26AWa0Zxq5I6nr6GZiysi3+sP
14FIOahTY14Plbsh1c5TG5Np0181ENpG7DHEzD2aU1V5sa7pNWC4GhBWjBp1WkFUyIb0x8ZtQRWL
XfmMCjCzciyk0YPQAXuqMpVC39sH2OMj/fNhJ2xmMbZRoEeamVASF04tA9jyTLOvfRajE7sZ1BsE
XjTrrEX4FhwhmqDhB3hwEy7CbpKlhTrCC3QwoHERjG9i6eFphGPvdykJzMeChx3aWApCQPZLJIqJ
i++58dRj/bnnFWm5QiOslnQX14bnRGC0LNEj6CNgBCN2zmjt6t17CM57xECRWKEN3zwoqJL7cmto
cDcWNVcP0hjSksfjPxhWZnDIAtDi8j5N2OO/CK+8sqV9Jsnk6cVqKFoVwiMCbmIvARH5uUX5Si/k
fKVP/pz728ai+C1B6XMTxrDugSrzDLXGjk8JM4pTx7t+LSc/QSqvAldw+tF1fwx+JyfQMsrAyRh3
uQjd6KWpzNlmN6VvDZVrMQG78j4borkUK3h2crmaDSJlCWoi3VYTpqvfiTfdzdHdIKOHvLvY10hx
cpR+CuvUkNdFqK0QGS8MwuILTBDtVkHGEi7j8ih4s9/OxFk6IUEQWszBG3LmEyFftUBeQ8aIq2ao
1I09RZXvKNcpGPRMYZKcbEK1nFaHTlRZNOdaYrEbc9eQq7ALPBdPCTqR9XGTuDfm9QzKJG35A/jd
WZJ+USjrfN50U5Qnrc4ezDHPZGVl85wRFEdCw9UQK5RZ+/QHyJksAW9YKcbHXspkJDHsYWwKMiFw
75yt7IHCSIwM30D/pgaw0NGdkdUgLAdp7Y8E8bhYVCE/g2+miKMuVvg6raskkBPDSak7yFwjFewr
E7cbDDlrR8B/Twh6//MwIcwHtL7eQNTHWV/85xKWsJLylAVzDZIHX8WpIzb9Kb6s16fuhB45TBq7
zVWnE+mGcJVjjVAgYqN2AlUUPJryflk+kyCuTcm0fACuD8PVUa/RFOIQHbl5kCnRRKwea2wAvruP
FKBKgjJRuPvJK6J9lW+7Z5StBs2j8sEsFuwJjbEzlp3NFd7On7wf6mLJbsdlPdo7qdRRLyGPLQQO
yKuZt8pQ3dB8q8rhJ2pTRKlt4zz6ALJuxPeUjLyuHr9hQqRuzjmoBvoxjYoecPPes3an1zsmV6Ja
TZiUxKW/2quDB6QXus5efeeuBuEklTlUAyhosuE1AS8p7b359vbt8pu0kYU8mTcHKrZ3syKA59Ec
2YGJE8l/ppNkGzTdRxn299h+I9LC58D5XEikrh8q87ZbVNs5tAeBuql/REIr3baB8qXgFqjsIUiB
eEILybLuu8LlPTV0C/pFPzz05qbs61EryfUstc7oJtqrGozzcUhzQdyEv7PswTYg8Sr7ZACXHYle
re23yMloObBqtS6QViPpzoI9iW7cFLYcxV+0O/jLiZ1M87MuOjVRV9l6GIPsWAohqNQYrSCDozvL
yN7m2EOIE2vrKaGuZ92Zvs55lN3T8IRp7Bn8BT/dvfsoY1e4c7KT2f5hfnydd4NlZ7QWofaZDNTu
fCdtjGMbtA3//UiVF/mqSMkyxhJY6f1VenqxDNJgBWkOSbjd5XmlhtCvAtHRfRPV4+OEm+9iVsgB
x38Rhxd+i9xNOG6j9lLB6oDfCHJ5shRQMfeyQLWgJ8uuHnXUe7kQJdHq3cFY1TftL7UnezypXkxq
dXWd1gtmpPIk0pBAc5p+TZpaTGufrAdq4UnFJKEK090PNUNWMbm1uQXZkTiXjsHJCwYA7c4+a2Qc
WiImzqIks77qlI0c1kPOWVBFSh2oGsVDLjcmHxfict8pt19VeDJ6ymxIGdPkMZJFTFAFTJ4pHr4h
Ixz6SPnvjIp1I689HUM+/loXCNIyYqsUnoLJ5zrOIJZewlJlNn/9Jff94e3dV/tKN8FbGZCNGR2v
NLJA2HOITKQNU1cTjM/nK3ZfVN7fGKJDEGtbaL0zDmhSpk0kHBk+NJQDtNzdK7z4YY0j1Oo+eALp
Z+qdNpnVKG76Ip6FC93Ch/v71lo9HEteay70Fz3SL0wLy7n7PiIm307gGvSINTnJwzI9QcKTye3t
pL1mgM9GpOexGLMeRDcZxvu4nArwwJ7R10N6RSE7DcpqcBI1EVkhLAesgGdtXwR4ErGBqJ2Vf3Lx
ldfKDPhia6th7jQ7VhwX0ASwYgwpqNHg6fNV0CzaSl+MoJVKkJGrTHT+426v+UumQcV4FUihJ0XZ
EIoPxVi+yGFfupoRdhfOwVRUTtQS+j/J3Cic8gOiWvNjHjpafPL89Zv/+hKVeVtv/YnLVo/3PQ+Y
PBVEZn3lB0vGN3Kqo9aQK+rySrGrApJ4TWP/BbiK0vS2QDjTvud1sr399qlKwjPKY5te2QV9yvy+
zYsb60k7sQv+nLQjDc8OoGvkcVWmKOvbyqbtaEcXQ0MP6LwXiw7HmqWyyI9LszcnI33fTh8eY/+y
v27o71kR4nWpSZhx+r1PWeZ4FoMhVpT7SSy0sbqQANCOR25xmZIscz60Koa4DUql/WKhkpqXnRvY
21rF7j6rUFR06kPUVaexGVnv8mXIbs50X0u86Y6bm1xu+MPvFUgwekLQxsgZ9+OchNqXN44SUcLM
tPodQo1KHRy+PGd7GZCPL67VBQOZ/oTAwqUT9GFN4YSSgIcNHrK41yDywyfWWy4quxxFKxnWFQ7i
//AGfgZhJUpqImr169DhByCksk8E7AsqmJ6Doe0jlJU1bP6gN4AR2n9NM5PpT4ZFHm8aDdft+dqi
cfCoO7paTkYd4ss29jFlrwkyEmYFlnXHaEnlKvNYLJYh5yxtBHvKTaweiOy8t8qOzS3uudbbPjrY
LmGcEd62OVroP32HWkcfUXP4QbVguHNBNhtSUv12hpR5HbPBZUxG2Qg/2KxZvvdaPrJ0R09XJD1H
9DDV/++3gxvq38AUqtVjYTVkY2zo8hxI1QFRban76Qf/cS9AQnOvRwg/his4tkMRXcEuQWxKH5IX
9UBsqBL4SPQBibfdI8uAWv775k/d8g1tLGYS87I8/HU5fo+qnolGo6GF+ewR1MShPf+bvdKJLasP
tbFZcv3TXt2P3ZtwlZTKcqGDejIUyJ7Kvb5HMBC8RTvGmT45PeqahCX30Ylxc1BS5n+DVTj2Kejp
mjShLgL74mbjcm0R9ghOsZsdUzUVpznZXUuMK6HINKfiN3EFNV2Mw7JAnac+M0GkO88CQLqTc+1l
fmC/IO6M7hTIhCoRrArulZ9fN8wa2ADY0sATEOKh9N1DgbW3jz/Z256TRKM0pNIwC/gnCrJ13Yth
aninxUmFw/5HwfhP3oh9kjd0+PNtQyfjjSv7LEx6Qm5Zoqhus1LPXT+CG+FoZnH2gOzDR+gV9R+v
W9j0vhl/y/u5HMSXTUvy67y1pXD5h29HPhDAYajNXl1PqvJqJDmAYyI5g6AFhfOcetEBcGhTXaGw
Cuv5Z3AyUexBjyXHa2ga7BFAEmPL3BGHCe9G4C8FKAoE4NxxfUyYpZwcPc60KeSejCywvwpH9rbA
7IDWehkIZhWqiW0BV2e3w24RUWUJ6vVj25UCv48/ptFf6rtidZOckhmKvcE60pEd39Uve6HCKQm8
uoTqYhjhujQH6+RIyUOjG+oS5EKOM1NIvHzAdD74ooegucZxYIwUwcWKP5GKzsG1UgWmxeGNQIzk
b0VdGFtwGlqCJeVFvB6Gbn/4O40YgCBlTspiAgHfrzntb7RN0FTNhpNQTu3MEBCO3ZI5IQvuBlVF
Vrwu++kKOF3wElq6W/JM3zJFbT9e+Oe7ZaCNhf9gQ4Bf0o4z9xwANukg4wue3Si5QubzYUQfJBSb
fg9PvZwPvYi3fsIJfVnuJdyIZ+55zFW9PlbzMGkEbby6KRJRFVzfS/KtKiK5zWkoBgvYXcFcUKBV
cUWVFheV57Bk/JR+QbJb4+74rpUsMruX4brnAnUOLNWBrolV3o0kDV26EiVobwqB5as1Fx/rPb+Q
2RZyiuXXwO+CDHxw0rRN2TNf+iQJ7jHnmsSSn31JFjoAOBAU5BcDorNJSDVOqgur6fQO0ai+VrgG
q0BqxPkApxwYWFiwHIznPaQtOlLQKv2Lt8e1YVbshyyjS5CoE4/8GaHVSbyIRVblxLhq+gh1wT2O
WFJCJOyaWkgund1k7dtYirw7v7ig7mbTrlqipY7wHt73cmIVEaIuvgJfAyiikMkBPJ/Bb9J9CGt2
Zs1J85VA/pA9rWF9Ygm6MBQZq/jBSDM9tTPC8z5j7omjkbfVOCnphkaCqFUET1+8srlgohoN41so
0jc4elaqwY6qIOF8z8XPndUPUxZGw75yT2u0l1M0CEHqyh4LO3cIzruyuGk8YnmIe06WyyVu5bT4
ARBRGlr2cXfSGayIx3M0awxGLhhYWZr2JxOIo7fCWox04EEtR3mOr4YLKxFBt8NpCgUAH+4JGjMe
crNt/HhJqm2HoS22bq3qSBgRqG8jBlpn3/dCe6qdAypYrXAtgljsytP5tov8JtPiiIgdrNUvNvxX
yrZvb7bxdoSTD76b/VLHQdNxxsPEEmyGPPcCPHoLDdC8OiwiTKZM5Eh4eb2vnxoFwmLFx+pa10Nz
Nsky2BC/OzVdx2TJ/7rZC5Qx6akbF9V+cvD2ZAyjvtcorp9W0Kuwg8JHMtF9I2+b0TyfJ09Z9u/u
6hL3FIaCfc1EoxWwGWv2lFZ4cjXNTLhH1kdqkFL1fb0piDImE+UVq8e43LVQiH82E+TH+ri+U0Sg
0r68YWp9Fh5OMutgg1dCvD+2c8kPR4zEPYZeFXtletF8uaZ995dYSyCNuqcCN82nMyMja95Xn+X1
Q22PJy7W44502ZCatuj0Iooy2S3GEN6X8BN+2WuAEfna+IY5WqtiiLhd4vWJ5PSNVoKRlKrdgeHN
UCkT2mll3N5gyKYyIq+eD5/ZNXKupuK9N7cd5OyGlV5aoD5lNb48Uznw6o4WRTU0j7/u9Dz0BJzN
QEdwHDIERTCE2fQkfBVGs8PY2vusm+bimTF3wKGJ1fEs/+5o7RoDPilZIn/8tA5asF3TGJlGa5P1
+dmuKwLTualI20XtBLep5vR5viFHao6JMsc+Ok0wkcskF/3mmrSHif1uSh2Ra+U16m3Pt8bl4TCS
2F6coLudKNN5JR66qEbUfkoODPSTwl+NpZbIIAk2v7/vrloQplI3ecUMeRqqLPDUVrRmutltoyiq
QZzLpncXA8Iuk0eIEnV8xFaoK8sHWcedAsomQyRoIYyg3rpZkB1KUwrLmxlyqfK/8HGPbJIQ8vWE
m5oPX6u969W1shP052d+oH25JXWCPimZ3s34YljSGTv6hJpJhPB9E+9f0PZ6R1lwCxB87m9XsFrL
SF/A9uIDa8yhpQ35KTZv+3j4rnMw0lOp1tcoPrtN649OfBQAOW8XkG7JLQt7WtqwXoI+bLGCZgTZ
6sekRx3K+GNOXIieyNd8KXjcW6VWRuHkssLFfuOHbgFEM8ZrS+ThHhHTiKVmPs6cS6V2eFt+L5n8
kcanl7hoV3Ji0+VAjxjpW+hDAOMTyf3agWOVSI+6qgFbApGLkYemGDQOGlC15BJ1aVZS3Mfs2iwL
ec/naftlHZRwTkh314lyLHaWDtSNc1HwjB6SlYvgGmq3yDfGvFV3Fyq76Cr7mtQW3pNc88ImVkdb
lZa8XPjrZK5BfahbWSHPzQ28T9ICcnBV8lLLjsvs4T2bkulNA9y21y0fxNo7Mf2B/gAXvSeOFIN9
eHkX0iADH+f77caJqbuLf2YI5jbtdjr2Eb5ZcnQFZvelWsFcDx9hDyGb1ffVicucCS7o9dIE9fhk
KtMSfDN+srTXyjTEe4sAJvjamPrs+sBi3hcFngXokFU4vm6AM6RqJtaBdLYBqrXZQ8gP6sOLyC8N
6xQL37YykMeOyzgI0KU7gYGgOE4IOHjZDIU2lzqkcjyLunmcZfSnojbDVEzfK+pXp3Dj5kVc/PAD
ogG5HNdIbuUid/ZOCNq7u2qKryBKZmjbLjhHSxKwaZ+/o1ksz+/rdYOSkhFJWpUT1Mz+vWmR+4Et
EkDcpsycTvRIOl9ZYfJr5elaUTORkVCHlP/y5JLsUwOyLvWWI1bGP1boG7wAnk8SZIGqNisSXO3a
u2VBNO5Xv+hAsjtDxUuV112zzmujtFse/bFxMxN4ikZqjHt61fBsCxEpeFTCv4RqbZx4p10uNDnK
skN3qzeUL0WlsplqBh0F6LyhA2mG2c09ARrKsmke7J3vrjm2yQjYhoBPPY4vYD3P4DjACDVss0zi
5mNGelm74gfN3szr2mwRJKtV7fqGKUfMd2vCRaj5ZmE45/xnEbQbposusOB9P8vZp3I/uW3akP+k
2seLDkj2K9/7jmX5DZD7dNbpbjA+t/EvS39kv+3YUbRPBNr3fZWfAIRMoSC/sRxKRLezez5UEDyz
PTZOYYwtfjEG3F8Ps+SH5sv1jMdD/TliMZTRS8jOS9HstVTzvXPpFQvecbP9YnomKQzYy3ch1ngG
nRT7p+/HxO++Ll/fjNmuyngQjcgN8CAVMhG7/QaW1kZrsvUJckKN/CkHoQpjWlibsnAPEbFFu04s
AnFPCQMQQklDG6TWHaRkQpeau0EWU/iEu0iW1XLc+f2IqxWhXIqySz58AlVJi89iSa5AIqHUJ/1/
bR8jYS5bh7uB9L2YKGjySWzlqBg4iCr+dXGnEYzaQdGXEfgREzqtSeqltjaRvdqmTlbxKr+OF1sU
dLSvFht3edwwhmx/6bSUJeXbFNuKrVWwW7FBjQudArAZYC/JontynxfbPm8F0IxM9/fFuuELem4X
4tcg/2blpJS8m285aLH11icM+MS7QV/jBZbw67fJJRVC2nV2hoXS3ai5Efqz7pGFXbCweMXqDqMZ
j3Jqdlj7OUWOrERwaalwNu2uRKDa9g9WjMg9wAI2IyNsfY97KpHuglXxyK88YzXFsde8Wsr5bcoO
cGzQdlzOi/u/ndkMu+5ZBKFbqoz67qlMIhj2U4Quzj2KHlrhsoFM+Ym2stEp4p6VFIbfktWErIhr
ltAqBvWdDVgU7ZeDAEUXM8bf1F7Tlg5tGk3CU9eq0uqxWtnz5sHHksPUF0hfO6B4vYAxCybONQDd
0KOJz6ujJyLF5KO/6pbHf3KePlAVCWMT0b6/3A9aqKRmMWBp7PRb7CPMu7/IeddwyYg8/q0AiF6p
Cg6X+N9tVDCzpo8vAeRp11FKC+sIMR/JsLABFqTWJDIVmEp7kOY60AWvZW9yl7AaFv1bZChTBMg8
VUxsmg7ELUxzlqIcHXpc1/2pRl7FUxw37dJqqto6pOnax7uRn9yshUjetzQl290NVHwlQ0gyRVw0
6oRKG/rjQBVrO3eOip+pdBXZuYfdA10VCJPqEnM+O8Jf/vvz//gRHMP71XUnO9UC02XOGS+8vmwe
mxk49qCTOJiHe5GoQ+JXOnL+FJ3KjQvHZ61SztHPzBrNj/DL2eineRCnZg2jU1x+EEwxo4N0uw2r
1DYRoFCs729g+4pKj+kbje60TUfjS0OFRrsBjvx6mUrImCC6yGu1FQ8poBaYlUVQJ31OKqV6EkW7
YX667S9cHwdtK+dxvSX5eUva4xGbHcorRRWQUasuKuEKGTJP9Fw29RLOC2IITxdFu026CoSNpHsL
BQhkFY1tnwCtWh9TSKZ4BahUyw00ieWR7Aan1p9i9dzgPC4HWJD1H8Fje10OQ5GDRBizk/Ir/Cbl
P1gFCSTNWt7TfJ/OOeWK/zYWZRJ7ZpXWz6CMoc1rxaMvb7UBIHgvohhg8IcLhyhvQZ00RI+dc49R
4TUUii2MIjMdAe5skRBi1CLKHs7d7eqDqq0JmOym6E1o5j6C30GOi488sa0ACgRedf7hchy3UJhJ
SJrwzyVHILxgFbPdcuTjwuJXRk9Gj99tUf36oLq6XL6x1/EGuwcfF621nDZCwS5TyAPpy6SV2BG9
PhMRzZHQVnYdo3R1Tme/FvMoREtjWeIwGFdS5PmJYvMHaI1VHys+YQjlC3DIX53kBh+I28GTdgYF
HwMn0z64BdPENNmAEq4Agt9xZ8sJRbgtGAoxJ8y3ZlTx6N01r1/rSxs0J/HYQGMCv5G7yit3gzEZ
CJmF0zKSt/fZNNk1F7jiU8OVqltD/uXpoSCToU3ItLfYXWg1fo2VVioDW0l7/sQegcXG79IZvbAc
XpKu8qOKMwwKbZOwdVysThVEdt306lnNa0aOCZcpr37IOWAay2d/nljkdrLpy9mJMjdRf7ek1jB4
5mGx7MylBaKCGEUvckCOXtLY7dXQrmwB1gXKsyyu4o3iye3OhFAZL3eS7q0Kyvw0LeuZJNL+w7kA
jMWdMPQzVerhlg9e8RDR1RoAFkZz38QYRij3nkzHjNBgcow=
`pragma protect end_protected
