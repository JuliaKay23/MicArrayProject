// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
c+vpE/SzhYUPn8UwUfsIO3WvHweKTanv7KOhrElhZTfndFB36sWjEnua3WdDEARmNpFMPp46NWro
IFJEim44C96l/ZAXvnxUShurdGObaF9r8PUonF4HxoOhqIomsq709fXVICfjKpx0fa6gF0ZXcmV+
mFrXZnk4ER7PWMYzmDnJKiAdx4aNlTWwmk6BQblgrqUpzIib+sFlNk4jbv6cHMfy0srhNYg9m3ny
cMBcpFjGeZyxne8L9Di6Ov2pdeNVIo178NU7qWo5qtRqknUTkg24P+u/7X7AWeYnEZhoTcxP/yaa
x63zElq3duUhxZwFFKhgMTWcd3Dm9eXIUZcrWg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 3024)
HJOrKe+8emUlhCtf84P8XVje3KXV0ffs0V96qdpI8fonphaXEBQRyq50ed0nRG283Oo9lfv2tbeR
2Te+YS6OGxpFimHsKz+JZd5t85QvSoElNn2hvSjF36CgRikt/VYoFqy4HttJkQvfdZuhow37iBxG
7cSqe90M/m1x3C/lwi9MSX+ZOFuA6D7eEZ6RcpWNEjKU1P8eDIL1YiXa/HLoDlxOpDhuWwVVl/mJ
L/uuEDDH6iUnTL++JUE+fF3g5jR7mjuaFT2/nIkFwBXYa88dhR8D+dNeC4om1HRCRYiSj8aAAgAu
yWlmE+lrcz2bw8k9PgkrFHiw9w1nMfgH8ed/VPu5o99CAh13c9lnyw7uij5WC+9CQZPFf5gI+Avs
sHZFQ1fr5Lqe7up1sioInUxpj35mcqqHS/273gdGA5IWtnUYktNi7kSjUuZjmzwNc8kD9fY662oN
Zw/GdqskYAxfL2LwtGDKQJceIP9dmJnrwGCkth44pD7QyKDz8/6mRDZeeRsBl+r7di5ZapK08Mj3
BUJ6BehIwIrkRvB3AmKoC51ePVDMcgEGxkURrCZv0Ilw8bJDghwMi1h+uDXL6hMPQgKlQqW5FVTb
S4+EAgjVJ0lzSmTTiHg206tmntMkduSb4cbuV1DfBLNrHp5Zia50jtMquL5oiJyC9PiV/4nT1JhS
2HoPcjYNkW7p18ApzfuT8eu+bFtOc19OCYFF5+0NWOXHFwq5jj2zCo0mQlqrqf3Uv9dYO6AKJZo9
9aauS07AG90soL+7KCggokXbVe1WxJ7BrXqNJICBsFLE+IwXKGGqPuef9xTM7zteuI7fIK0oQP6+
78yvVLHpCa6q+80qO7wcuWD2xTsOn5EXJ54d+zLDrW3MN30gIaVZ8pZszHTuR8h0mxpaZ2NKAJ8D
rVsd6RQMDnLMA+nr61FCAukhL6SIgaofMUQlgTohn7FpNF8TadZm94N9SvKh6UxPbAdJlojc8qj/
lvPDORZt+4UZQniab31OcjedDm/K19e+iWXVAmL5sCZUTLWd2P+yYmcIQr1WW3XxEVulMA7AcSid
0cjvyJWaAzGLXfZp+UOl9ZSVKK7tCigcWWzUZxvb0lLkkzAz19NKGeek4PR1ISnGXmestvM9h4zd
DZa30klBOYviPBlCukNRNB4oEaUy3XPODiORqYihLwVzwHg5GvVYAR7eL9SXX86Wt+NT22BIpfxh
Lf3BbaOpU7l/hqBe7D+Sdzob7DFKlCZyg6z6rv1Hby9VGShItAk1flh6Co811hNzYxYaTc9ExdZm
0Et1qaDvkbpycgcRVXWKsc5fxtsDth9n0cBBeEVxRfXfesu7DCun1HWlQg+yDF7/vMGjnrC4/wuo
uOG/BgDXgGPAavstrxi0KhWK1Xa51L2S8qeovmhLsqPdRMatY61XnaXpSDss2D+1CusLs/cVDKEF
9sqVFFotJadsSvA1giGRvAp0lc9yAO7UdaWxUPpezJSFAU7jM8SuOgPHQa6ypeUsyyWpNIYEmeMy
dXMUk96KRMiKdJRK6j+kAd7LL+wJ7mInl6INtCZc6Oi2IJeAhU+qdSimifGQCu5biW7Nr1/a3A15
NNG0pp6VuV1pIWRXPJKb7WSp+oBlZuu4bxsI7U9MuHx2WzcjEjs/LwQCJO6s2/zJB/UGByH+RQl3
ma7r6UQCwkkC2M01/MyC2C89zidTu95rUC7dPoLcBGVxLRn9wrIjvRDZfLaIXCtaylt6D3JmU2I1
tjYxMUI+8iuIjMw4WQ0CbtdTGSHeFx9mQiqVB8ihefpKZHo/nIROkiiYsL5Fc940yV8C5ca6R33B
0xjDeXmuIU9HkT4KQAVuTxQJpizQeXqYwQr31pJn6Cunf/Qg8uM0PyurcpQMBDu22CAIysGlPNGN
Mr94sfZ2sP2VbHv4QaP08tUIfDun5MR4GsoOBdNo6AG+5/jBTEsM5V3PSjT17BnscRsI10IM7ocO
zh1fSngfyuZBLy6GBz5lqtIjrWw2QtL9KMHty/L0VF8GG8Ny/H2jMcQFy0g5znaXHTg2IH43TjHk
TiV75MC+K+O1JT5JBL/1i2zkgG1J2lfH4RYNR/sQxayf16BLNpbwIy/kbRH1cr0pjpiK5FzY1w6K
unchugzV/DsDzN6iYH2fC0RTmsUNCbRNPybSyTjPjQZCl+p0saSqPv9HpASWJvJjetM9e4XKJA3d
XQ30FenT/Ht7u4b4zm1B4EYqj9Pl3DoZRBqLvOa6H5FGJKYZgl0tYEKCx0RiuCA8CZwHcXelJwD4
YOk2yRsc4jBFUETKhAaol0Xn9eghYFETPXmT5PUZBO9+1SFN5PWmSlgWK6MVWypefDUHGheiS/vF
3q8M/ze6yinWDTfK5Jy9xjwixv44mViQjXBABx7tb/quLkavZdczreqDBkjOqJ0ZZk+iqx9ZJhH6
0/ps8RRyL/EAB193EHKQgroaQ6osZ9ZGESfbx2bpkWCTnpl/nwotabFnLXmDmf8Pr0oq2g8iMdy4
P/ykKGndj01rFTVZepmoitfOnoGAtdp1KI1otzW0+6pWoVrO7MA8dbwBaeOCr+qlGqq4cMqvh5OH
AAvSj7wobMh7nWWYbu3dH/DF+01p9KkKEhCvBFYTMOOfPYqzJvAdMWZR5AcH31/n+KXke6Zww/SY
zGf3Kgz7oBD6FYfsgXVDo+PFxh6EXKrZzOFwBN6xoxWMHRk9brYElexRl/minAX5CEF6MCG+gJhE
5hLoc50Iu+jXLdhMzzYfrCGRhxJOc0fXl+iK6nFe8MV7JzB4vrpUYcNfWcmvv9+zcFF06FTLD9kS
vQ45w55uwc1YirZOOxOGirwKWz3xZ9MkAjqsgbNvM4VQOx77k/ZLz7ISmtXS4qqyXlqRVg1WxTW6
yFTUZDUfg3ZRtejxBiUPb97A+adhphwaJeN1xXzSd6ILtaJwkPOSJeFe2HdPh4brU5q7qPIJrZzg
U4aUBxJFlerd3zxUHAOBpbm+eaU5J+/wfI4G/m7m1g2ovgtxmXPHSkS8XY76KkgEkUXHKNzdEFCy
EkyhK+IoettOrDj1qXNDva6dowlEh2zXNxqlJD+XHKtCwfyqRDOESL00OxwjB0umCj+C1G+mnDeN
TUoNAqSq/qamtelQ5kaPPDwBz1NaMakdcJmQrAZsZHLNf327NNgL9xjO1pjWEZry/hBpKWPPhZQw
ZOKfEyL7uqcrRiAkTDD1IaGoRTbTMz9J79QhGvU03rTifUdHPAlZHzt4IHlrHwlkZWC9qcwCtJAe
0VXRY+HNgu66oe6sHQHfTOCB8usplyzdvHy/79QGXLVqz0Us3igy01dght4Hg/krvBZKErmKJmiR
as2l+/Ept0O5AVzBLsvUEwrorCxnVHJzN2hensheL8F1tsfUaMy+15vaNyHae2XLBGzQ6tILC8OZ
Kn0DAtzgf2ktne/rwj8QMoA6d44drKIeRwc+XtTnWcdW34fvXPPEBjSL1ehqziqzJRjgk1vrj7VP
xjTHPEq6F5cgOV9nZJY7pmNrU5zHte6k6wM/Q11/s6AYY0dEyvQQuh04yyr1/GW9qDNohn3GMepI
uPTHtkiR6hL/cWTv60JyP9E6ZownGi4ZQhmB+gqM5zVpk4SuzChHUMEx8wqE585BG+hjxXiRbznv
Rp6jdEzt8u4kQ1G3pdj7R/gS5hlec3SQzsoSGY2SxA+zPJrWRgke0UFURvYtXElSI6okgPzmg5j+
88Ib8UYsOBt26mgtD6FUCVUH/E396Ff9fBiRT/y4Ow47Hyhms3hxOddC6f6mhgZH09bRrnPuCWW7
4gqQ/Dp89wr2lv18mvOtkKIbrB5GCMHJ2deqNRT4b6ywmnVecGuREn3+Odhrt5TmhIQTruc5yj9i
mFGagpGNORBtrDTfLzfTdZB0VQ46YQI42W0yXYB0sebmpVBWg9ZP4HNZ0vNmWtMBl01XArFd0r4+
755bblY/gV077ZNsSVY6P6mDpQ/L2cEf/7wH622G7iVzJVsaANggO77mZQPhxCbthm80rCJzUyY/
addR
`pragma protect end_protected
