// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
EPWplE3462qUsHVUA65xLty/+YpOh1iBt7Ootj1YmwRbA7Meh+lcAx/5nlQRuLH5OikJ+Idt6OLj
ssADqPbz4bMvCxCrLJQrtVwlIKu2Jpa8kIkqiTnil5SN9KZGZzkT5o2u8PhguGa1Y8MaOAQo6ZP6
Z8XhphUctfC1m0wldGFGpPB4SWcA5nGqhSTuwbCzVZsQT2MD+tOy32TY4NUoVuNqIkrak62WycoT
lmeyDasuOKO9ikKbw1hZOUSb3YctG0eGPqxtqS/r9Hllyh4pUhgCxn4rLKQyrVzpGBrHDBVQW+vI
t7jTyswnrPeS8+nMKMwlcQOf4EfSH7/TRvUEUw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 21216)
o+qQo6SfNcXSVzExD73n0/+yq1OWJjxvSMRwe77cyi85ahLHGedFPcy6W/YG3zCmpzFD80WJm3n0
/NXltBMVmkC2u89UQxVPfptVgBrnihks6uVSUnDK5pHnLvfKqbynJmhZjN04dwqXxxWzISO67AtA
rD4InnShYp8OXWYqshvWtRp2Sf4tjbAUYP/Umi0x/guG6mCJRXnc9QljYlfIaXjmngu1O2gjG/Yo
PR0MuR69tntuuTz38sWARKzGa+wJqr1A4MSEOBPhSJ1LtyLql2KjV/yPuwZ4ff5I5SRhFlUQ8IWJ
XkMikobzj2CVQolgWXs74gIEyY2NXSpFlfWu6FOZKFPvmdwNw52+hGTn9IWPl6bEUd5AconPWP1V
edr2Ug9rt4irV7fcDJ8NqGfYufOarz7a+cAMs/6NXVpZeGlrSYgvD/DizM/dS0YxSrgcWaxY1K11
+ScHXGW+iwxnJTrictEejo8v+3dRBe1vtXFE5LCfzYKfJJzjcuOQEutDjOpgv3BAz/GWiSXZF5Oe
EomGYcWPbTu+88BIVAP7nNpOHdKmkd44mUaH2p07pvUNX7E9SpWuzWlzeftqW0PxqWpL0av/RldC
jaUPbywMEdHeRe9KmmkqC4cUGb109/1GUkGUqNlnhyKXxsnFhar43trmmOTdfOMJdeVbG//6iLVD
rDYRUNzkne1Stwj+aTL0EcaF/rIu6aBV7QU+mHFiUDthxirTb8x3r9q5sFbJFR20Or5HkOX37SC2
hLSsDrYTlGbp7NLx7vdAB1wbVVCvd47JAZzHrUTxzR9Al0SXWUA1g+kzfqW8hvFQpFw5JwlrEdQT
5j6QRb6toax9FbDH/70mLsoOm2917/ILGpATUuy1G+e4ISySV8w/rKBvMoxsoi7euuZIYAAI8OgZ
sjXf35NtH6V/vlQLYmYDlpJKtNZhISdDoJ27ACarpCSR/fHpeA8it+RFK+ISwhiWTDW/FsyRwmsM
l8ZHuibCGnMT1IqbWR4Dp+vGLi3xSDuVAM6nOiGFMHFyp2SpwaXNguCpHhtYrvDLvWRqU3QsF+0R
kaipf3N2pHvdLAHF3Dd0XysZYil+o8QQxbR3v1Th5BQwuG3+vSTR7WV+XbZPlIYDRoNCxcCmiUhi
maR3gwieZHwogxAsx6i82r0qcHjnV8CvHa5v4EfPmuou9+yttOAOCOefGGEqC6KwHl+akXF8OrQs
T0wOz38L+OAMuR63WBoZl69SmkgRo8U1r8S5iWkp/PHnKF7Aj9ZwvYEnc9+TLBWAx4flFFatg1I6
NLGJf9QSfmhfKRrhbuRrmrvnSFd+x5vHF85X0FEp7ELRiR1rhqcoNcg2bk0oCoVHA6kXEvpnQ6oT
7bR41avBbwxfYj2rPctTWxDhEwklrgCbgMPrNfAp64vN17vpP+1l0PIiwXChqb2TmYWxyJ3sYEbz
8zAT2l+fP0QP7loRuey0S9h3nc3adrFfujSXNvKMyHP6ysWAT8T2bu3Du86arZogi+Mi7q7iLZvK
AZpx7vy+4aQ59Vw19CBIqbz7BadMsVnff95IcIyocxwM3Mw7Hx4xEHtwSdtT7GOsrp+oWqb+W4pM
bnf7fvsGL7fiLeTAfWRY79oJacNT7TIB3LTvpRaDp0Cgevw9eMByVUigSlhz3nRQqTcb5WFaYw8T
wmT/LWXGI8iOaSm+0G1fnt0nz6bbYcIt/GPS1qvas+MJZr9pY7UDXiPb0Wy8yX5ia6QxCA0oMbH0
qk/ig9mXUS3WxyQuahlRLysBN1n12nYbY32vouE8tBOF4KOlRsg7490sosk3FgcUotjyu818wf/B
/eeXOk+vIpUAdJd3+JpjhWDZ4lQY6YixU1p07DH4TGiT0Qtq0WLOMdt3c5qI7iP62+47pH8qu7I9
0q6BZow9yLejElLRmRBm4YMp8v0Y1TKzDqfRQgxMWAxiJscBO3fVb82c3d7FfZ6rkbvlIC9/ADAZ
cEGl5r3OO6GTrhrGFvnGsk+cMyq1crN7berRewiHzbCm5fU3A1PWgN0Nf0MtRswv4tvfIfrfzjDI
kSSXubkHt9q7yb+jBIv4ljDJTbJdcD6QUKPWCF6kRELQsdr8+wmYE8ztRJB42mYlA8TTovvUzkO8
/8dctcUAH9GF6aZqYoT1wRT1TyraKuR7i9/BCx/qy+KHVw9OVDdBVIMyIdXg0Bv+Ja96muqWMzx9
vD4gaV/6ah358FNVSNI9PXDufCUvulDmeUo9sN9DClCavPO6R0/pZYApv6nARO9XrtRXs5TWmjIy
UygU0T0gcGQTBEfxShM/4CXeNT5KK8kvH6OlflcMyybcKxhaFY6JR0Hn0gX+dgAxiWH+DdBaOMAt
pnizxsA9/fAgg3YGwvbVTnsYi9h5Y62Iy8gzK2vwI8ycoLNfjKHXvaYww7qvyxmiWGI5mE1H3L1x
u0aEb9kkifI02rYNtcUfZc6fjAEXhHlV8xTdoNdsbSnik/iDJ9NbR/MK8k2HI2k4sG5kW74dszzj
dBhI0fga8vo91TzVQuqVbJxrrarhxU2NbiuZKDOk8//l6kKZ5lHfLexkIKaot1lLPOW87UvTthYn
RwfQgstQNIMjPf6QseZBtEKUcjIXrxhzmBH8cO0ZtERDuLMnDerZr51QxcQu6p/ejO+eQU1qU2jN
9DUqDFuRZVXGsJfhWjtsMUThulaOraE9/i3x4idrog0JyCiTcogfH29gyNg2xzEfYWXfzq1sHJ5/
4HSDa6slqxeI5ZwM4L4cP5S3ADoDgQJWEEHKazxCF/TBwmiCqZ6d76FmYo7wlCo5Mcc4RMXB7jvc
XapUKxCOWHuXf9CXrqmB69KfXTMcbpcpUYcmbtK1QDSdpwoKmNiTYn3u3RGWR0QDyMXc8D6q2/aS
C7EacErTov00Yt6QHfu78Grm4S9vgbHL6ZZ8cngYterzN7le/PJG50Y6SSwed3QZMWjJn774lLci
b3nq8M/9qDx6Uuws1LYfwOhMuFlShrRxfyFC4dS2DPAqJBIwhHoksZOqAEXSVuILqeHuLXQuBHjq
DypN0dKKtXe16sH2BGjno4A+kqJXncgeVSYTxp0xROOOgIRevNe9j4j3N7x07G6ghBDAdBAO8Voc
zumfFkn7PuZd9wlqzBKaLll/Qthr5ojLnbY1njwAjhAXmt8+R9BQiHqNDiYt4lz7/ZXWzH7DnG+Q
ktopVdnISDsZfK2ExNcrIDDgJdrsfeoAJiwIuHgol2algnD1O2imB7PPzEbWQY1tJRePVpyW5Py/
qOlBozR6BBCXbAJH5sKJExfwd8YHJAU1uACCFRwu8Q1bgzGtVfYyel28BHgYGnOZAjXquUuGJLg0
lIjH7tCyUeFa2sv2p2fn6UWKOKKaWTvd45G4dnb2SW+yetxJnZXRntYCZqAcx9Zow+2y4qp6bZaB
IcfoQy9QddUKdAdcAeiS2Fd1SQgv3c7k1eL1XoSXwa9pyr+v1zor7tmKkZ0ikr0/Mej+8+jh5K+t
rG4kGuNoHJZQo9KYKn3cCg1J9a0BHykc577/leZTRb6EwD2aVyn4agVFAK6QgV1La6OK4MV5Hk6T
Yra6Zu1H51QkUzHF4om9yOjrTTp+JS2BvPggTKWM0nWKWaK/dHe6B1lRdITf2XqevgGnKl7yVqek
rjnl3dNFHTK9g8NojgcUyWqGcRwXCfN1I1LKOoWXHb64kzwlX/T5UBpaULWLTT1GE5iI3BMhr/xr
9a/RTFOtIRs4+yDqOxQjTHYWyTthvn+n2gr+GHCgZDZ/lW5SGTG3qo9Ns/6Jxl+5VXwKR8r17hHT
JSv5VTSVSEmr/OsOKLgiGC9+mml8HnLuIuZ58ZV4ktKIzmI45Cf2vlwFHo6CUjIuPVPl6q0tMbpZ
cScdQwNCG9tuOhmsIl/selzd69Wuls9z+aMHFwFULOW9OxFP5a1KOS5SUscb276K5RE6uglCZjg0
4big1jaJC9vVFc899oMyzxTZD16KmeXjRETz3oqCPSBblSxVZ6Pe84AhgdWCavC/Rm70UqcaP2ph
LqEcXoz5PcnflQ0SvV1YcM2mF4yocU9T6AaicTZPbArhVcyjQ1I1xym8UiwpYWD2hVeZ0X+Npb90
DqFRUaSr6jsBpJU/dxqeN0ZYstya277sjuJs+DpeByJBOSmlh+COsaK6Bc4MRUPvazZkCrHNUe2s
b8IDaGiHySAyuXrHKgGF81DIB8ZjeoKen5ffWfPJ4k9u4JJQ6S7S7jXZ6S3paZw4koL4VhTKkAY4
JRNKLZFyDtyGQ2c9CEEogjxugTf6W711ZtVg0vSWwOa7VTcGZJamtMsBiEzL4PAgtvZEF8PxkcmX
Mz38eGJcJTMoCs6nqmbON2zY+qqqt+vOTCFD3IbsUxVbsKaCgHMK0zTGxKd472Q0QRe10FTKW8Ut
k4tBCk/iyEOrAp9E72kBJwBo7L0z2NzfctD6eNMKsHQPAd/GbL5LilX4Lb0bA8UoWIup1SFIKOam
i6LWSxy9FIGR+5jD6ToT8EupV0W/jLRYmbv6mCq4u7qp6TdHOCtRGa8319EHZovJS+JY2SZ59G0j
BsEylA63jOJzoNUt9V2MMpGjZvp6LjXEJGdmiRpHXRWGUwLlLmgRxwUdPPFkVJe+XTOtoJThlFcj
Rg/lTaUeQCOJt5Pe6quRo7Y2k8AzQcet9JH9m/1/8hZigB+zLQ7AVMueNrnP4ofq80acxNmGzQ1i
GlNUSnYZglaGh56/jKDGhLgTOUYWUFTlYoc3/j+3vE0akiQgE04r5VN0tEcoNOmo7yofZvS56kwe
MbVkoLQ9IWlbCIOooa/0r8BA/CUnFE846Vs+X1n6wBlaKLFB0OAMXNg3eUgqf4rhGEKwnr44cj+N
VVnfq/74VCyLkVs2RhIaptdgCcP4XFEORSzRnBbhYKM9cVt5YaBViaQLCEVQiJW3cxyNP+yk7+Ck
pEaokCJYRhKnm0FYQWyubMErTFXMlPcOT2vXILvx6sd9ymycvG6P21z6AbjEAc2VKTHhLct3NgiC
s3QjWwGpOe41NUUKqxGpyuohjpt5ge+yAmXjCazI8BN1K4daHpa7Rmb78w+9MT2xrHK43lwxas16
dvHiL81iLNmCYsLcoQaXji0oXo3LqWPM8Sd7iSDQU7JlIZb1Xt3Mg6LnA2Tu3Fobd1x6KFsvKyy7
Aaf+ETDvnHIXSpE0kiY2PZ3WwtxO0uEq/1HmGZeP+QBGqYDyQxBqJXjy2Wis43xdsQtPT82PqZSN
9k4qryLWPHMGYGT2Gj5PhMKc3AWI83pbr6hap9VI73xSeF2ENsaZHsJwQLVZpgfpBkrTy/uneA7s
MufWSGCsU+XWdz6U9xQlB4aVbURNgU5asqF3oU0CWvqB/DxBsfvPM7hx0TOuyX7xIAeRG4d3E6VR
d0t2ci2L79/lTGgaH0x/fx30ao/nufBuHycCRj8Z2NxHFk/JeM0dAV8N7Wo5NU1+RLFBu57FWI58
NihhFKsHD4ozLWQxQtVljUtt+LctLr5RdKMI31UeW7a9CStckU/chXGzFHsDBWv7GVm4kjzWLVGY
2u3c5pFhK7WAEOZxzk1yF+MMuFMzVM/c7p5hnQIMmFESNkNtFlJlEgFfPq9TXMtMYNTgAiPvtGzA
8uWeJL+/yoN3oJ+n5EQEEKOj9pSe9jQdAbbb8969bxMQIgJgQ84SJQKSF07cDescILhx60TRPEy5
Zr1ZV0pYoQbCccrE7tOh6ysEdI2z8RgunAv910e73sW5atw76C5OOjUz0y1SRN7wevws7qRQEzjx
2iiDAJrRMfkV4I2yHOD7xo+L+s4zNQFz2n5ep3Dc79K8P3zKFrN0vW0ToXZCXwtXQifqMRBxraxQ
+MQG7cpA2oa5lapBad2yCNq7vhIOiWIx1xa/H4EkDGxdsGZFgYsnrBYi/4HmoG12gPpBLPYSieMk
1zuedjJcmjpg2AggCs3VY0lX7QlA5wgHqWH2Vuv/tNvbIFpF2ZnqDxM+tCdhZVFjz1TLoi46XpMd
CahDAXbwEQkkWTQB2/XTq5UaOZeC6fxuPwcLW/YVPfynouwxfcVaXtkiFTb/4k/qGfBInRs9nIsv
cvroEFpjXCwocE5DuzVrnsV2s/KwDa067UwrOMsvbuOds1DEu3r41adsADj6/by4A8qeEzABgnMZ
irbESWrlEboJTE93xgW6ZiEZ6OsWelNAp4s9OAxmdYWPxlwC5wJ+iOTVJT/VIFuL2Z/mhA+IvqPw
+vY844Bf8grjVmqMfiBWJtkdMrHTe1K2HkF44MDFh9NgLtCJhno7deJGjkJmpqYSZGojxwGk5t7q
HfH41/ulBp8koPl9gzbADMi3vMldhppbr6JcqXR/SdU6DCmbqy1lbV+Sl65x/tDP4Qu0Fxonzmku
4fY8XatDOnzgXB8htp018pVxor8XMCuEqNw1ZIPSrrDX2N5TEhmfhT4TJZUxQqeAahRgcq5LpZiE
uZk6V1t5juH5iswboK1nIE+QHYPl3tQ5xDz6Lz1SJ81w01kQSrSehg3gBOEH8W+Fjl9/vTeqki4Q
ml0O+/9wD+jy1H1v4P0jI1IcOwkouuz1klXzqipjhNMwbnabt8XpP5IpgrzNLBl5mnIEOrZta18a
FQZDc7zJta/r2rjzPbchhQdgyeSQhG2an5MvZ+47DKWkfFUQpbG4OdlvsXuarsI+62rYg+Q2OI3t
zwsBptQbfbThDyJ1Dr6ZN9SeeFh3BmU8dbpDxrXyeuEIvVeZvOyvir0DLTImBl/+RWk6fxe2sgE+
IjLKQhfd13JUg8LmD1y5k360MTvnhgM7K+UAf/gFdeA+P4dPO/b2RSXXk2PPH+iKOc3/gRuR93yw
s9wdeAzgHeVuGvJxga8+kLcSqfwfdU8PxY2JNgMGK/rZNwVjJ9vptD6BGLqEHUs+be1k7EpnNBcI
V+CxJ4ICNi1Ij2KCS+ffEEXPBqMbPk//fakUDYu8csmRAHIP5eIZVxD44fiNIZmSNUTp25xYyntr
Rhe20JeFgHMaMFzR89nSz9iUyw5MT2cLYczWj6XoSqs6R5Rx85WoA2cn2tdywZgL8DtnK42FPgLr
WZWllFq114miarI+C3FBZQp8V3v8mGh1C9D9c/6vAIOR+95jYTFKLXnvgjbG8mWCYVt6SQhWgWMm
znR3qvIpz8kEkxEm/o8hbRtRmv9iBDcbxK+bESk1R0Wg+Y2yMoAmd8ZAe1ysvBTt1iwglAc/SnJo
rTH2eZagZmOR1GMOVXVfmqRIyB5Ing4qyyxuPhp8Zfe7PThvDgof61nhcOqbSvROXEMJ+DC0Yig3
AQE+V2LUaTf+0rw2xXMjHDt1lqBlCpNuJf8fBY+j6Vq2pXuDsI/nyoGVGVaA7T4cMp/oQTQ1PiPY
TLFiGyBk1oZBa4qp2nu1SEEbpmOuqJuFn91Ci+SVqVvpuDxAD9mR4xfHZ2Y0kVTb6hfnzU+CKUqm
cDt6e7TdXaCTgg3gHrGIr0GupaBClWTOg5KUVo/n+cxkTPEv0bOEPn3f+ud5QICJhSuceXWYZ1cC
rh1jkGZCfx7uEZUlJW4D10tcl2hnEekIwzgsIZntxLF1tR+y7rwUMAHFPuCx+Tg+Szdi7Fy79kBR
+FG9NtbPXGsIUS+rMLtXMuFnoGw9A7u14nF8TWQyJhXaI9sVF8bG3cWUdzPjRQyXS4dLP2hU+UQl
NIZJC0TRYqfKXxRFk3LIpZEJ9EAw9zZCST77h9WUWtwXhbJ8Ij9Pu0YjHlUpuCzYQVSBymMeonX/
BlnFZPERtXIqdLyMg9w9DgtyUTO0tZETnslZP8Hc6fgQh9licqmZ9nBY5xcEzoNiBB+J/z4Ufn9z
Jq1n9oyyn+XnDEwH8uugqXi/lY7zuu69Jd32khQmwGEIB8XKY5a59ClatlVR92PYp7deIG5gkOC6
YCjT2rNnXkKos16yGOAKcdg4j0aqY5TJsKjGA9MQNyWvnmwZn3OXP0cvEtpqZ5MtrABZMRHM4RRJ
6yGl7kAMTWhgDPMS242E6W2cMsRLI6cLx+6m5CFBo1YzW6j8u8L22VxdRJb2Klwt5msxsrSUi9K6
/hLZ4+JoKhTHTsWF5Z+u4iKCg3hecAMn09x4WSjz9XfB3eJ22Jlb5cjpw4RHVwtTNGi+RF3jIvwv
U9isMb8rVhbgBRVaJpeO/Apo3PkXFGj95fs/fxTZTYG0VXXY0SUWZS1GI++X0Bv8r2tgWAkfm24Y
WG+V8Ju/gObMEWnu7UFZxfI+gAfMDPxSPdhx8PmfwVJfqlHCTxgMXHfno4Q88nWtCckn5x3lY7pB
IOeNuxNR65zg4HexzO8j7OSP4yNS7rjEbTeOmIzgXU5lVU58rpOIY0nJMUWhLO55wEfXMyJ3HCiv
sEktQpUA7spOpCF+lOT1wOWaa+WBLLvZ9IX9ENCOFAM06noAYa10Ag7Qjlg+u6kVGY8aw5gVppOf
VfwxHjbNSDNYGuKIBVUZKVEovFc0GQhRSdKKQTRj95wdLiK6x1ZZcJ8A5YIzni+0yrXkzXiZ2uOm
jZLXO9Ej096fY5J3RAWzBwHIAaZf/ew7Fw1tOUAUYXa6TO7WHcnFkw7hOpr4Weqibz+Q5bKzYOMw
8XDovOCufNyJeNG/0/ptn2OjTOkNxZqxTdlu1qAmR7O64fYPtrVeg1lW25uuEDOoj5OnOhqkQT7H
IUbpN4rJvI88UE+A7P/gvw5+XnefwPv2QHq6/zcW0w9w65U72djuMQ6tAm/dsIVIaJhthqT+enQp
0zVOhyqTHHA4ekD2egiaNmn4p5D/ptA0AHp22nTKgaHlggUhu/nRmwh4MwP7ZhaG56dmGD5w0MJO
qCVB+BTnstUmwllzBzaqVN4oJ8+qQubkkEAdCaPW5jiOjaL057pieT/AWogSnhYd+EcwWHzpIlpw
1mHpodlJaL+pOFUv+HClDUhtiMKA2yhzSHxpkg81dq4KwJogG2SobBeG2V0unLVEQOLHobNoUXOk
APFlPze69gfk4iY+DlDnwN/P/q/PAeAjcU5ZBRFKWbYSxh3gTYR8R18B06mOKKP6EJy23vu0BCcC
LMiwXpgwkMl4n9QVtx4zEqOHFOoC2lUWf8sYsofCSwqonNhcw/X5lIaI7jjOHPBNriWSikUVVz+O
ow5zM4h46wAhTxV/PVvsbGd0T72FwWVQfrP6bqMJwCsJ1Td1/HGo9e0WvfDh7N47P4QVH5tAX8wj
8lqW/x3+vErC/0rGLcCblPakbCuEPemP/TU2Zuv7Hw6i0LYHlDR8ASecQHX03SW8GZnKuYnyPTbj
cQd+MpyeJz/KMHfjkSE6HcY8eh3NCrYzsMISp95BMtWqFwazEb4rrrMtAV+Wvgyp89ciYXr6MWC+
qe4WB/fMPzx+wbSJzoNqY9G7xo69yDyEOzcx6uCfVFAbAOqKsB/lD20w4Fruop0Fl4Ahb5G6pSrC
KCnAiT6VZrVnRe+UpQuJuK3Idh42oPd2d7kf9NRaHgDfbChmi/3XFz2UxCnz+2GxrJBoxM9G8tVD
KU2enD+mKZlD2YFgf4nvN6V/rwNXG1nEo8sJl2DAg8oLUJuf7stYGuf/vSgoxUfR6CYjOXA9UdHW
Grkvi5NRMLWk6NV5UMrwubfSAgTUmcrwqNpv/a4OYZeyzE92sVYXuH2Wu9lfMOR5r0QHTTPOjloH
IqxfPNFrfXwSLniHxzWh7Xj8odh0pJOyz4h23bXsOnRA75M7i4GvPz2PBFyQl5Ocb+tu46/LTPN1
D7Pco8cCgT4RNrCosu4LFzAQHh1+cXCo4+h80rmgkYGqY4oRUtwDkCAFXUYT8KgnnrUHvec6t1iL
37kHonLWDnbP9DS0UPES1hZ2Pp2ZThAnRjKaH0iL8VwhnhDvsm0L8rD0sYzE2dNYKcbCGCfzFXjO
Yxgi5jHhLnmav8qJdp5gZNVOWs+n2RWo2OTGnu+MQfzZR7UV7W1Tcbn1MmgENyVK0wlzxMd/8hWT
9ekk8ZSUbLLCkva8f4mSnA9suGotlf5dkwGyOvzduGLtNgutAzNnlfL6KttnPVfauxqG5kHVvOs4
9y5JxvObv8mgN0ScfrmA3q8+oFLBQ9/eSjLX5hBcTnxdzGn727ua0r8eRhErCCncuNABjeO74NTp
QDLZr+HhhtrSzdNdLLkMfazTQQShm7cCBGTsKLBgMCrS7nlo3ny/LtEKsPb9XYoCqxdgEMuHzZPW
BKw0saPc+me0TA+PEfJD5tGQ/X/8BomOD1p3wDmmudHZY43boXj2Ip/5lCj2lVhOtNeJ7KOcNYQY
u74VemNAAxKjSQ/tvn1+GiW4XRba2lI6zLCu8RHXG9SlbQdObA3PBtIzSPxgs7dNPJHYJM41cxsp
4r+6yv8UVcvK3871TS6VaNctWmjeeRQmOXy2INBWDDzZfzNF5bZ6IsnYZyy3e9fxyLawQCj5ee96
ZFoEZWX7vh28AQ5iIipZSdXvdfgirZ7+1rSYBboZJ4QEtIWPgVZ2OgwgqIh0PmO19k7h+4F5+OMS
m4G1PHCD+LlzDsHXWXnXsqw7BEd5Oif2LKy1KBvaJqkocx8ihDbhNunojAVA6PX6BBui8kmSj1Z/
U+CDSO0xxZS9QvLOC6P+myyLTGR67lj4rGDjQJTidFtL5SozpwAMd/rxg2jN9XBxLRuHjx8rGOqu
VCJlrHQBpD66yJZ2++MIYw+IPyN6LoHrKnzisXH6/DUxem3bCS4ICfhChspvGW/nuP/4Jj3CxIMI
BFuon18MexlHEuLyBBaeRjdUX6o21Sd8lOkPy8Ha8fayFIsMl7DtsYIUtF2HAoL3ZQjSGrLO8coN
v8pYBH5CQjidpsKdYxaU8llBRfql/upJPi4ZsJZU0oy2nN29FHBrf0/TR6sfylETYi6eHU+Zx0Tx
BNxMC41VtAiCOp0zL4mObmDoG9dO2VaDFomSWcIl7Xu6+k6QC7RtWCt03Z+1+HSckjauxr+smMbF
rZUHUTFjjZoe1Zuzm5LOytLvKkmSSlEwDP9WlSo69OPtEmayX9U8rTNqdZxLpncu5OSp2MJiiUjQ
TUJwqqbSrIZ/lg9zHYc7KqIrolYbXEnILLf9rKr0bexFyfzqA9j1jc/P8HMqMcKSVwaIduKpqDx1
xtViDHOIwIAJV69B6n+VXZ62OXzSF66+I1WREi2lFZQfsA5OIxM8YFzxjkbjrIWa8s8rX+hpp/I2
lySsjhajNvfZNV6YhBbqaZ9PZP/RNlfO2HKgd85bEIwEk1v+Dl8r+H8nMlw5qPdBt+nuRMw4VVaG
J70GYcYpC0nzDWgSRfhbTbduRvyXte7kQ3mTTZD6U6ZSM2wVx6psyU2QqH7slJTvJe2PAuoApqm6
XLGULD9Wh3q83x8BnvT4oAKmGsVjQD7/FM/5CpquyhHUxZCx6pGrXeYXNCFLJCEXq1pksViOWtG0
eHyOi4EsUpWHEwRG0tc/yV3cHjIxVm3gYy8Gn73hs4CHdiOg+rD9zl9lNb5Zcveur7dEhj1JOQQ5
wyB82wPBUQ8tOocr7Kb3w/Zi/67/Wkh0Ay3JprBLoG7YA3JMLuWhjnjwAh+CNPw387CDg/z4zGqE
lWmocspVE2IKAVJu52LwPyftJivyTNlJOtPtuGEELH1aazFJHFt7pKutAbeVRUBD9omU7KlJ8cbS
2vCZLWNxpxez4kTYcKJCT9SlviVWAhknODterzpwABOwpg4UfgwB2TkOePxm4l/S1shxwJhN62s1
rkdWA9fqmQANPvQQnI2CBIb56669Q4oC+qwUfQSNpX87t2rLqp+9zd4WhKx1UFgAu+AHo2zBIy6V
8K9MGoJqD3qc7R7yuMJhqvZwdwBepgbcoHu9aHKpP0sd2OdIc9OQp7jmBKfVrqQiXUrVffcdW191
e9jXM8WlGIvLZqMOgRjxQCQIsUFBsfb4JNxcb0Y9laEkO5QUde/+gT1zNNFA6fdr/5KGwiIpBH//
39lqW89Zvv797S/H0ZfRHw1FtGFToqbpwSdU1Q0Fk1I9hcRJFFZX3OauGfhfPfLhI6Ea4Eh9JvEm
2ovVAHpjYP0BJ/Tmq6I6E5uFDwn5hvYG6qOiajB7dnb4XjtQPqy4URSlewNKNYjToNwLfMu+vBXC
lYlk+tSngM3KWmlvni+klK1r3oPClTfkRRCBazQzqpxWGWihnnSC+RgEWx5ZgSLI10xeVk8BaGA/
0Fuf82cqYzKBy0x6LWCBQkBmtLrJ/PvT1w536Emv7EWMChxBvyPAjT7sjmY/82cc+dy9+sN4N9gc
wDyGOFKx5SM5N6o5woM3sgzKACrIzlHlW17sZJc5RgRH22QmAdYXdIGqJGA3SEpgdS2S0BXsm9tK
5xSiI9RQKT85WSU3I5Gamy2K1Z9WAXO+xA3CtcdWhGtzEYfLQVwGZdKojnauHG/EChuAhS/Z+3eJ
sELzaN11i6fzf1GRLd8+794fLFu13qML4kNgDMbR3ARQVfeY5o0vbXgjj3xUOn1FG5hbaS+uLLiv
FItkA5HCUuvQpQOP4aFVYHVeewwRKQK++dTLbGndz9nHTZEitXDMAX8HSkJC4IPL1t2eAabNmKTe
Oxc8FKEZMxGMP8B9NgPMdssrUa3cP/Lui/yZ0aGhWzr9fyhzRZpyJKL0oJKXzSHx3v3XxpynLK+I
HEgbT6ZYlrHIeJX6zEhoHkZI7+msTtUDRuUBrIcCmrbnoppYir6d8HGYfaBHg/+yd8Cht8sNtfdi
Rv3Sa3rqAUiAa6D+7f1ZK1pYCy9dC7aUh4RfCmT7S9KXNgLj4xiGWH6KVRSRRkKddxHGafAAmafd
MXnMD1+5FpmNRJHEZ7OGyfdFDMKeGoIxalF0wtB0I/GA11vU0C5HRQknveZBb9RXHXYg/7gOGncg
whRnmo/V8EnNRroZbYGWudO9zTy+pzlNTXif5IcmrFtOlTHz2LIXQSly5SMECmf/ieaOUw4LU7r+
/HKhBtYCqTAu1KCyVT0VL02BQs5MDtcu3UywLOxFa9ClrBsqqNnBKW6qhzIujI3QwLryzQ4MzzWc
vTWwDCyrUCHbYvdfdq29w2QEsfyTgwFP+uGjL9pt73LbKrKzYMG21e/Qll+GnGxTyXRaPc5NOsRq
bCP49Suu+ZIYGVuwrJBdB0nt+FIlK3vosKYR4kpra1iQC7f1er6ledCvwkL362wwxVyeYRDGKS4b
1cif936YZI20q5emlmh1noe6EdwgAlQL3vA42q/SsHlMeJi2uptVWjigxAxTAB8BLO+ErUcWNSCJ
nnJViG2P0fI1QIJ2jC59FMDUqG6e0+V6WGOd7j4VD7wdH+3Pph9nGr4GzpDc29aSlrWIsIuYvO9m
LvA6puF9XVVkjvQEJ7quIZxAYjljUMd/poXh5xAUIFdOktmukXGsrOqE0qc4J8Qicc3HFSneU3NW
wX/ZQTNRd2RPBCpWw5AKCRnjBRrjj8xwu9/fjK/eTRkpRWJayqC7jfPpsUDmLKiZ8TsSa1A5isuS
aAnLI6TvLTC0wgpmCdN+1z155p/nAoZrXBv6ZSZy0Pku+0YIJ3QXta9tU/C9Q0R5cQvruMJw6PHW
yaMP3moI9GGwzft6AtzgKGndTpHKMjsoySf936MIxBa8/KYYrZajeikzPQYBl+kdhvjdLoktVMQR
HCmvNYwXqIJhXcgCUR9UbYkmDxq0E/lUpO8uGwOMUU9PBDaOWBRPWQACW4/0FBQt3URB7BHn7afX
gO15eEZfAf0GokDrSwDqhHYtD6YDEA1IZ35t3KS0wIhpnCZ0vVOGoJCQbStNB3qeVLrRHboPc2rO
XInVHzfyYwoM2dscYo3ZamCku/j10t1i1neIeJ0a3bUJGMc/bbw+jKLJJo/Cu6iaY+JeymVajbVq
YjFoQuy80mY1aaIlfnYoWALF1I1FYkVZuFep1c4mnCWAajxpazo8JdY84L4Lao6yaYxsBKcXoliZ
aXRZbY5Sk5nqxlsBCdd5nuMZHEG02+aVfbxglRFKcpDFG9zlzu3r66B3a8+vjiap7e9sEFpuGwA6
TRzfsE1YsfS0ILSC68nM64XPWLm7xOAtO3sAcsUub1hScsSa8ack0za2cmKICnTiupKLDToo6CX/
vUoXIZA1j32LhC2Ex5OamfaZpsixHiUN8HwKvsBrn4a8f0B970iSssZILzQOvdMbhmIhysH7nC+d
COO7jLWiryNjoN3MRQuacgEL/L7KHlrIoewQBHQKKEPOC9kZ6/A6L6ONylOCDYNfwOfxR5v/4Qa8
PDP8iD1WlV0T1ll0COGuD3LOQ2lOw07kmu1cNQw5JOvcTVnum5xBlPixoN3IoWQjRd0H9EN+wf9V
MNJ9SIsnN6PY+yP6zrDUyH0BwBO1IrOO6vbKQn+jad3qJ5Oco5dyegonQUupQY30CHTEIcKXnQRf
ZnsobskcJK0sQUB3Yw27NB95if+TMYiUscZ6zjFfmsubUSiX8nHKaIuQlJMclfIbttbxsEpwrQHN
a+CR4Obpzem1X3vCtj5qXGP6kvUMynT31U2T63XT9NI0bs7GNsPWxmAhyervgHgtIKac3L/n51KJ
Y6JyTjA7MA1sJzge6lPkO47qfkyHvg/0wko3YbIUgQNxYdVfGFFa76LSxU//B03LnCMIwuEczCSW
7kCCpNFgcXw4L3uh1gIaHIctDjcm903kjm6Df+YGOYdKrU29cgR4kpFKTkY4ZBKksoeRZBZqcam+
iEA14FK6Xq9dRavC6z0k1DsILB5rWgao4FcnQcJlOVKAN5E64eYCfPxno0oCOXhcCM4PCja/XIJT
jJ5t1v3D70r55NqJLBIjzEJvypTz4RrQ6u8dfAN6kgCfhuK7CEHkAqcAo5ufUGRUhSS4jPEpJesD
lekuu52M9RN53r+9YrT98Jk3gOEnxtXS8M90u+3gIGtGQpiGHQguBs1gec91AozzMr2yfiqr9Jf7
MW0ZyAambEZGDrUb9b1uvzvcQcdJdh+dBPqM0EpWF4Cfy436uB1QF4EReE0GQPL22e6o0OOs6QU1
jA1Fr+DYkujon+buUkHdSsIcgwSMMmH99OBpYT7AzTzT0Y5LtFSBNGxgUcQXJ+uPH1Y8wx2M7dbr
PkibonHAGJf9XHXSh/HWwzYAjBzI/Sv3MPbIi+B/nMEtKObZr3A23y8L1uKPeV1OT3lUrNEnP/At
u9Mb5DrpIPh2oANEOTKeNfElp6JywBMgQ1x+aPg1bte0mjuaqiBbkmMi69TiXc5iTtfK6uJJDWgF
PrZQrIp+Yku4+psNxdy1Fa6NM4GnyYodzXA6M2mBgg+CuS8AJn+NEGMeEmtn/JiA00vzKubSB31G
/+ZP73xDn2ddOKakd9opA6NRv7Bl5VkVJs1x0Z1ZZS/OsPZ5Lm6yzvwe6ntEZPqkVwy8DYakd0Y+
1TSDcOp1K+3xTfHldcEMXULPpFUBKol+/lnKcM+U/gRKo21PYeAbLGoxHD4SRPIWg9cteoZ+LyoN
K7ZGTlGtxzHTJh0lLAekVnsQsXz5dhWVQ3dJZapx83tEnkEOvuYsWZ7uq+nBj4nW90tEVuDr6AJt
dCWAk9KAgihxOpyCk89LjnbESgxl4CuvuTwtm6rTIfp/CoXvvwarvnaJBbhi6RnwU5EJ9tD79J4j
IvSnrxnpZgTXoEPdJh4F7Fd4M1Qe+8tHj3yBoEGfDgLv2PyM/x6Bi5ntv2vGmUtdlZwDHkmqLSUe
WzQZ9UWPL2ZFpDaSSTHkg42bJzmQIwi9aFPtPSyWUDULiHoMW8YzX611/lD+Ub/lgLDmrkPV5Sxz
a6hsyV7brASVStq+MjX+oesKAhDY8JN4rLXmt5zrVhkSEldFHyKMqmlSgBHU2VSEfm0a6uVgBf64
7Fvv+UbpytamohluzObB0CfeyKHEoFLZtB6/MQfGZxsl8VPM8Akw29N4NrQdjPYNl1dYqJssJeP1
o6cjRl+fJ6dR/Lte91jDxxlO6tKZrmkJdaKMatJTUCy42NAWu3XIsTDVETbdouWkNHXf/T0YRNOc
df/sk9vytcSNKLthhQkV0+sXm6RAh/4X5A5iJFOlrwYEQb0UAWeunxNPAoPbg/akTe6zgV8gcLZ3
yiGVLxCkuhV2APl2vzKpTP/G63JS1Q9Xn3lG2GyIrdyDnWET5N5OjwhwCtqcRV2mh7W9RetpSOXQ
kww/9YQzAk4Mfc309JtgYx+K8MQI9RPCcJngC/8CbHcQLc9a6xfTX7k4JBMbhihXMxfKd888Wi0p
KM4vxHGw6CWbBSYGB4z9hRaWrx6j4BDBUvsQUWK7JksTvw+P1ShhdbGIv9iINEekboGSwNMNIK9D
fHXRa715zYBAPL8p8HGqUzsg05rbNJi+4vhod6DN3LHwIo5CEo75R/lOwzg4N7yisVYMcNKF3jlX
GJU8wqnQj56F0Zj/MGgUDLDNnGMZzbaTaYuhvtvgiQroGcXBgkjRGViRs/PMNF9XO61gXrYURlew
JFPtRi87SPO6DYxmHtmbvC5bynNGyLnqCnTCxyEI3x2/b0U5drJCwmwOzFXKTSF0Xkf2fBocMcQq
8EAISqE9CrehGb9NW2QtiwOh4mN7ymc3AcxUPX5YB1VqzGEwl25VHbGZ1SxImbuwHciwQYm7Ukxy
4TzeVPw6fswwXa66kPRpEquu6/ePXTcS5PNHvAMrsnHCi3P9ihx2djUuaQiK9RMSuSYsTh+euUOl
Uaww2dN3ActXGfEGiYvYNVZk0+h0xio/2xLHvWsh90nBbUVAOBeQznL9B2orw48XhbMTXsUvFVTC
gQ0FrGXMKyWle2o4vPUSkVQ68LR2a6xu2JNRXzaU3ONBuAMuQ8YV4kC7fqlxwNepjD2KVZ5EHS11
/cqBhd+KnicuLdJu8DxVhYM9cua7SV1kNQHGTesv2D9GKymX37d9mgsjPRta7/IEkkhzfe3XfLIq
nVwACYV+TLNvDIOUhCni7rFOon17lO0LzFdXEwfCtSF4Q/YOimAazESij6npKH7TzFm8U8NPQXKi
iTlNExOBEhHulvnO3dh15avYDefAfUH5L1KNridNgpfxJjH4y8mDps0yJg9pi53CYxxK6+/eq9Kc
qPVKmiklIKrSFNlDatpE7uEfc2wsHVAOb4o33sL73aM9fQmDyCmfuOrPkgC85bJC0WV8UM9mQUmz
GkNdWceI4H/enVL9AI1L0cRvVhj+e/zYDt6CwbC2muoHSWBoCsA7zsDP1wPkgOasqUurirs91f5V
gsYgFitpE166gGrq57kcsbbQbQiY5LLQUvltzyg9fLzj3gUrL4dhFCdMcccgBpjmyzD6zAX9PIDn
bIIJ9LYIliXiYW9JEfuXnKzGV1gbKIUGfIxdBTtE2cw7fTSm21uQlouuNkSFZOBf/m6zgDWtD7sV
59qd3KXsjlzGFf3MxPANfROotphMk29danCIIalI8XveZOzAnkZEtfYqCgCdU6M7wFNYvq4/vn08
rVOyiPHdaRGakL2QfkwlFX+mtEyq5Ih6b5uOKh2GR52r+nndKPqExUVaSISousRI3je3bt/bXW+p
+fs4RFFVrrvpNpehdX8eM/995qgBEsqvHjRD61TVop91UN6ZIQchUaKw68/WSTRStewyXRiuwIgR
kuM6JagFi7QvPFK1xHeIati+mmbplVehepIHoISwjqsni0Mgto/ZBMUxHthNlkthBN75EfMeC00/
5n2t65eXPnTO7uns1F3nwDpC7M/+HG+Sdhc9ggeSGlzQxGpcGYFhqU52RFoZR4/rfEAzN7ZNuMs+
UtMqqucwjnmgvP3Xij5fvUkToFp38+vlrD/HWj08Hfa1AUPZdU9mlObOMLxcQ5Y/OBVE/26RztJS
ZM/fnvzJX7LbRWWHeq7Kg95NIohAqO+iW7yRKyziWUIg/OP7ldeLlPvi65TH/Sl8F7RsBK/3ph31
bJBmZl2XXiNsqukujNoX/l5hElo4ciwGe4IauIbN1gwQWfuWCrxhY248sJvc354c9TDM7vDhUGWV
M9H+k6MydVZc7B4AdPHlC8VCoKK2F1/556GpqU3GwvegrKWRe3v4MOMgE7+e4K1K8RfchAXxuJTw
WA+AzATCFbZuaStV9K6N1MYyjuY2f3urlUt9P+LohoE6NeTVXKmy6WAFC2bq4V6F3r90LC82Csob
9DSRVpDEnEI6ftWEsQquCjZMnJQi5Yw6n0CFgsrLa5Tp59i+mEgrN89UAteIpNSq34E4uNX23Ec4
kHWoVXYcIjTyQrxO0X7LzRoVG4li2K4olawg1HtVq+tuwXzrNEMGiy5PX9ZBgythhIs7RI+srcVP
9AVnHXZKAkH/LIEwTfjP2ihE1hFq4MFRRQzXaLWVELg8pcM7crLaJ9/udwLWF1Qc2/7vo/RGxAoC
FBqUH6k19iPmbbwlZrpVo53c7pJkMGGcUXyOqsesW2L1UUL1r4wP+OlS0f4Jn9fFPoqLBqfF0KXG
cuaQZ26g/OVWZKlisOAKVB/XSg1R+nZg/Bwr18PbnKZhoHUAvqF1hvPnjM90Ji4/zRDrIWatTwAn
TkxoHkEDWg4tRhPlW+VgU0DBsFFNRHJvO89yJGJVDKDZhDWWquX50BxNDiHdpQWUr5sPrwK/Gsbi
9sbzMMIYYloLW2dehSgVmnazpcqELRBLT4XD1KizAnxNVuTGJCREhQo5/uWzXzz64HWkAx6IePYq
Yn5pT6lejTGQb2wTDnVqs8Oxyw+/5pECOee/569l8FZ9j+fLpFzhLrKgVsM7TvXzgpdsjJGOeROp
wEspJ1ZSQYTbdI4+yNBLJZri0Vo4xfTLq+JZRYTind9C7kv9Z/UqYItaNQeuv8sCwrMBFzh3c7dM
xr0aibqablIxZOcyBdycRafJN5cDOUkyJ/vQPigpnfimybBV7be23gvUxk03WyA8ULmuB4ZV3yfQ
laFCJgekU20X66SSpgfdV+ogAPKwDeZwp+6vyJ0wvUJouLWYgegsHbXHKm9GVZOWtEraEQjSpGlO
9PtKnfOdped65LVeE7sdANyN0AGYbcGdZA0aUZLnQjuOY67C5w8B+cbu8lhlQ85+lze4NevHerTp
zYX1DsKBR9+DaGPIj/pCsit0YkFBylfhA7Zx1Tj5wVOEVnd6OvnJ4VlmstqVXM+QdCt4bGrl9dhX
sI//nfXiw8mACi06uYzwnIHh0k8az4reFoVPXiJ6ZBWzF7W8EkkER4UabWO/NDtjVWEfyTSsa4b4
BXSJJzQyAlCxPgQEjxJn4yBZjYbD0xY5/VwHufIP8wRerWhOM5qJG2KIUmJ7nBD4dRKIpInyyZVw
ipdgbpkRTMuQEbcWaLMbl/3Eflejxd4UxzuPWolEToKzurSkkuPEeJtVfWP2pj4KkaDZ2spkkyN0
v59bVfbKY9ks2CUxEahNK+K1BTPM6Xq9T98Ti3agpJpuaPLqbwQvMNpg2l7unN828W5RyCuOJNUz
IpKMDk/r0/tqWbLTUFtJWtlWUlvejlG/LxJQCqtptuCcbDGOU2m/vlpPpwjszHE+usU+a423bRVh
Cn3HVTOpdcrkTRDgp4M290PKpI8cKENDRfL9lv6okJ8GLduhJ1RJizAMoJvX6O6qr1eAvX/82jRe
P4HpzxtP58rMVnQJDH2Y9BCYsDioMpZ14ARUStZLB4QHltg01pMWQIWfNoOkFuUxCXHah8JW6kMK
xHbKYeuXZc5MaovMvS/0cKHuyf5hfcKUIpkG/u8L3MWPFuHgqZUvEv8+xhUyaNUpo8bS6aE+UPg7
G1SHjg2GCw4hBfBOelQ1OaqvY3Tea9ieAfKzndNAiobtpxDhw0d8SiZRXgoFOPRod71ZcWAEEhxx
eRe0bdRp/XoYNJIWUMTSA5BjjR9opUpm5Ej9T1I1+VkGy6pRnWkdx46LPMJgsDu1Ir+3t7R7UBjt
W4yPpTP9LMbvYCRfaBuzeC+PJh3Lz4yVIiTdIXriOO5QnLMU7p9a31XUhoUeeDIEWNK5e7CoQZwQ
3E+ZmjLgYPgfEDhl2eiBlACKIQwwP9uMugjCndSD4eeaXwanbyXkvppdr29DcZdiDx2PlV2py7MH
FnsxlrFdBU1ov107HfX2srifLOhWt/zAZItXa56Cvz8hiK6XB5IYn4SVdcwI8/Br6NfHy9vFfp2d
CrmMfn7v/kE+YBMunF1fg9EgQidc9i7SjjrXJ/J5wtn3yT38V/NbhbxhMLSo5tI8fLXTnkA1Y9lg
P0nnYbua6vbV+z49R3pcwEzTCca1WNShvN8QkhobUQJwSM+gyI+oQ9hwXtbqY70+oRbQFLnRYeV/
7RrDCptB6PoySlo9/7q62Uex0sCeeNBrRtL+RK0ypj0NYQO5ejtP8eAJYhYTO4vwR+f0sk4P6m1J
a2Bd3+ABH/jh2WeMBXXFQdZk4xa9TDxaTytu1uw7k0YaTHskXPU2O7Jig0h4HU0sC3AZM4jAgK8K
HCwpO/W5W0XKcjhQo0jZE8dN3Ip1+26w82awgDFWsFwZfv6Rk2CW/yCVVRoYiNWZ0G3rKMeXjk/U
0ALOZtguVKVSt6b/+locZ4CDzNagqBnuxZaPMEsnxaovCNTy681w4iD0k5J4c0PkVLH/fC7wN7Yf
BlGzh7UoeGBuV0qmQ10MnPmT4N8ranbrVq162bQKk98OTnVtGrWTdYBBjDJU7gbBOk4DY/HOjzgh
sK5m8+oA8CLFWmWCBSsUklqR2U3pa166CTHf+Z5riFn3bxHLQtSSMqn8Ex8ZP60uZBcSeR5iSaqm
Qahiwcw33/hIvyyQpjXZPqhz29diigLULkl+XcxSgKIYEZPtKcOqKDxgIqmn0H7bNTDSpM8nJuQs
Au6WcuFph3GfrAn26C83z17SXNTOykwcNR/wbLqHUgxTrt4+Ua7Xw1g0UJ8y2Pt8nU4m3O/v8ofn
7lPoglnwhQiKOVRdwyn29mMTEfYCMx6YhuRDhmhYjZwU/bTKVToG7SBMPG975IvqPS2mt5Re/EY4
pEJf201C59t8MDpTl/ErAu6DCuYMi7iPEsRpZESHnGuxnAdx5qwJDoL7Dcv4IWKpy2JFbC81sj5/
QqfHsxNDSehe8QrQO9tMZ0BZZOHkWpGeOWFuQB+q9vTdd/9vtaguMVDzxeT5HzCJ2Eh7bKUyw8gs
NA1EMvggbX7WKRgyzEuR+E7hOJT+lMrlf9OPt5vma+oc/ooGblNWPp4jvR5+320JYPyfK91DwC74
uo62vL8/3SS9MwEZXYHOICWygUKaKRMz9BTzEEQONug5JhQWQUtR+ix/5hjx2cCGxNC+c8cbilr7
XPEeKz4cJCLp6vkP5BIxi+KHkubgibgBaVazuo0vu99ykVYOAUR98mhzLY1WsNa4Brt9Fdr12hsK
/pPVF+sUkg9ugQTWaLyyQatt25qg5Tpiehe71imJJ7KXPkMPjlPs3e8Aqof6r+0XZUJeoUv8sG+m
BQzaKl3/H8n+8SlthnwiFm442ScZ+Sdr7Ea7mi8+JdDBxm+GzIPyzmn2luyc2mVwtp06OBd3NUmO
01u9V0w9QvQCCjLSmMbI4Ni9wYd5ysQ87jtXxp685VCCtxv5Zey+S3fFpdd7dJM1XEKMq/6Tw1OE
NdJJsKnFrRsl0xau5AHvFPwG/gJfav5kM6Ngi4ex6qzG6vkEvHYqoUqqGD0cyYZ7ap0p1fRzuxIM
rnA3H7wbAMSFQX2Nl8QZI21Y19UcMyKDje+tr1Ev0Pdpxlh0cIE94xwoqlUA9aLUpqMOHvvvUSBJ
ZCVlnfYog+lewGX1q7fT4P9x5M0J7V/2xE0+DAQ+il6wX+xR1296gv+SMrr7bn8dnXLSPJz0b06Y
uQM11GnVuWzf+XRRx0XjYgs+RtWRmg/S0o2yf/FaJSQ4Rzg2CZQprPT2M63LpDxF2b6b+Os6Sf7h
Gu4nwaPNVtR+C/G410Q4oS3OQ3oNZ4dVQDiDlERD8mPdiwsOorx7wnFV5KiqzwzpBf5YKCONF+53
FtMoiv/JyTAHDmZX2gr1DaFAfX3Dqdudtgry4TrFHKmQDOLJXG+5gcQyIifIQ3GyssNezlRlDAKD
JWRmlAsDnHBan3rWOBlK1w3NoS1z8XaMuxj8HfTv+ViZnYUalT5s7qZmlZHS9tAmIEkPNmnb+jMa
dhxyb6kydTEw6SaS8ARZVKOQkwiCa6dttTEnX9I5YZNdqimczGZ5froKhR2OY1uux8rI0O3/Xlhc
CWlbSKXQX9+k73JktD8ty2M7S/hDcnI0Q8pEOGcAo6vYTm9Q68qZMwJu6szkwdvAjKkx9VJ87Bx6
TPlUtVBQ6rahiv1O8xMjhVjug10aDAZJil+T2EiEOiImKxy19y+H00UgOuPRnWC43YkGvKb5OPW4
fluz7bplCuow5oUCdrIP0J9Nt+2KBqRM6S7UWHh0EQqrRrO6RDLxF0CA4FEoVwms9uimsO/+4PEd
ZKD1BVOHFusz0n+1t5r89V/WzuJB4FDe0JmhOnGnRk6EbH0EvyU1zPxcS/2S3Envjq6Bl202RdWy
pJrkb4FC+EPJha2MIHRkTf0NNtL4kCONDZWvZxBlKNUhUCDnc8dmewd6y3TjFcMPO8CyZkscIWCL
ip5BJVghQ7UUe+mEm7u2z4kBcw7Dq0Dm8XRiQzj/kgHB6FXiQUBgH624i4emcQBelmNYuQFCN2Ue
uueGUZdqPaEvP74K/Mz6u3cjunfyDkRmKJwoHJdiyCX+xE5DYXIX+ikSwhKe9hP3NDRLtweOIofF
nKu4JTlSd7zg2XIamQoML2kbZb8pr4TeLjA1ODRJ1aCTMd5YVsXnLuKNHztiUBbF/D7JiEDXanqt
xIDNk54Hp5IjsxTxyae4Qx/tNbepNA1k4Fh65Fe1o9a4u/wLNKhvA5sqj1HdULV7x8PZJhnQxyTf
ktRz7JCP38mxeUwM8cUWAR3INrOD1f9dF4bdpJPzDXv1yVwNwhQQu18rD40YzP6U64XgmnB81AGn
Urq4/bN13rZgwH3vOzhZfHaXZ2Y8MihFUOXknw6j4jNtREkx7k10FhhBvPExMYj6fqmX7NqJZ92V
f9gRD7YM5X4VYVEiK7lttsKuhoLLVA32hdnGBJ+WXch6KzMvu9z0iZ5ySYQCpoxcKMS1vftfj6lz
SI0hq8+IGPAcUKs2+/ajIsmJwRmpslazb1Yq+FHoRw5Su1u6fdQB9mLsD9B+Ye/xbA0/hOJXV6Q7
2bUVavKunWvjvDnTCEMTB591RP0dFaLtrr6AAyV/pLtKpGUBbu6xpYimOgyBnVHuMFM8O0DkSYE+
0NT8ojQFqvUFR+PY8uiy3UGxIwIEH4St3pb6+T1IHVceX/7PcNs4ck83buArpkxZZyyaYbRyhTDS
GB9yuWQV8MGkRPJqL05qOEchRkf2QoxaJScg2L/38BHZS8unBfRhMgBV2hD8Q5Awj5Z8BILNS5+b
yv+2tqHj3NniqzPbxpL5gA+JP7xO+31nqNdbCht2mrg/mecIcyW7ZFYyrQ7YUYngXIi1NpDERkad
Smy0CTcqoxlWgbJYXjmpKVHw7dX81izAfXQp4Qehtilj86CWEFGGY9VtqUi/v1A2X141UZXCjaG5
M8tSOfU9RLQk5z81CCMjSyF8f4RufO8fvJQDwmDyamnaSuQbgaS6Sv1GVGRVTFTscNUxRyJ2MjzQ
lABySUt/dlBTy0kIeS55W7H1it3l61073Aklpfcx6axS4dROkkXfWBfOOgMDoZBd4au3Ejbr66Ky
COkiiJpTQ1CCshpOR1sp9YHDjRo7ijIavHVotWa4eqHLtSTfF4n4T5ha3RQ2BDQMEwTpqdaF+nYn
87NDo6f/ElQ0H59VergRskbBmO2mRMSk7vWf5xASGC0gY1rOAtbCizai+YVSLZj0bLn1u6UqLLsV
++GQ5cjEfRPy6B5nQPk/bB55j2D7w39LunBi3xUHANJ/8XFHna3lGQE6+4wyCNMPcoafB/prIFHf
tGdAOBWIOVFioCysD8PcTM30QYezqloZk0guKvWfd3glK3uMrN9D6kQtMEnFhfTipjcYbiYf//JH
xax4jov0Q6RNym0CDsGaLjT6K/xBQI29FjdKvwROQ/lovdNusStFJhs28yj7VMcSBwMuB7R4IrXI
JDUesdzEJ8yvJCewhEqhxKeKAJ5TIpQnrIxhXDKVj+7ZqulcR/hGOZKTxxasSC0VM6+WGd/mq83y
TpJkyKHJNAdcIndskJiDlFlRuM6QN+DzpoHhgAgp1GGc/b9lcl/gDSc59vzNKGQ6FgiuFMlPD9nt
KUD26yy+PfnjdkCBJuSe0KfzOla/eEZJmzh/Q25tDTNWUXYD0RVcsYmWtnRwwS4PH4GxTUFzJy4f
T8k6RI7Vn4BCM5XFNkoTZXlaL/llUs7t1C8X4V8ufjuF7ibd/ZzJ2HDG0eL+LjjNK78c59zHgnKa
0N+Onk+JOwGk2z5UqBI+rnyR/usiqtJpfkgcZj0mNaGm4sgBjx6d/YUKDisEElSBxOAknmLe9XMZ
bHduFPk/Yq/GeQVt+UzzcwUq05CqyA7nE2+f/3FoB6PKCvHIJ56oKFDTrXQfPQwagk3cjrsX0iO0
9BiRH1ZByvEB5h0vJb3Nxycq4Ni4DCqXfH6LGFpkKwUU75//G2lqjjfQWfwkx9Vsni3dGTz+A4Nh
xZ0b5s0Q2Di+sm3qT5pNyeXpil4eCvXqRoZlJkPb6VJSfTof5KYzcPZHm6pdHLkD5dVeBzj3qFLq
kh1lNt9+8p9/05wF0zzqOtfM1wtZucnIXw1yI0toss4l2s6xlk2Ldffkp5uK0AhFljsBsH/6/3xd
A32t8XMC8iTR50C4cd6Sk2dmb+ynhNJ/4MSYeO9Pa2/eoLxK8lmy9pTxdZNWPqY02gMsCRDUT/du
O6JCB7z1ayLsIL4reXg+9wINiCAjt2WKCOqRLMSKiam7UfYAl8XuwaJ9mOP8oOtqN+gKuaJbv+OT
4S38L6VNMbkszsOuC2F4+Z3PmTyVZeXDZm1QXMqnpTtUbDACDfqDUUbnRPgcTX1IBy0OllySxZ3O
OgW5th9OtWT0joR9O9WRYOUlDB7zHE6IYcy3zL5U6xiK+c7TzN3Tv5KK4S7QTZHNGEanFIaxlIfl
rVa/IgVEvYWpmdVI2QMFTFqcO9Xhku6YS3BYOArF0vnziFWT7zITUGzwBB4Wl6zhPU9dTcGan4ci
/IWEhsgEp6L1H+11W4rQFAMBndY/6SoXhsa7/5cuXC90PhL8aZ99+wY9CkWh9l1Ot/YUKYlOk/uv
WLPT/TeUmT+exmLJ28bcXXpErE83xpzy67gTIYvRedRCk6JHYeh6Plgb378HDguZagJCd7qwVVAI
A1Ugyk2JsiMOndZwZmbLTdJeSQgOM5GNeS02ah8kITQjdNpOYhiINO2nqiYMbx1reM9TSz/dP4Vy
1AxOMNYRSqgzgOGyCmJA08QT/ZG/xoRKJTaCyfuV41BS4GbhKCH43lAqULs8njurdHmGGtFEmq8e
xnjoeV79FZ7Xj9TmjmHqdv/OaNPMr70SoLbknPrkdFje3xndOPShLdEgPWgWf9tjp7K54pAG6p2a
a5pLU9PHrjJn3sqZzNuV6X26gehIess6uu6zLj1OWwdIic+dOrQhOQHEo41Oda9wSQ2CHQLUkMPf
bquuGlIbmjsYUQ28SpJogZoKWyCwaqkcqbykMrli/kX2K434DgUOKTv8jtOkx0Psr6ls9TWCL56B
0bdaoifLV9SJ4WACrbHqlcNYlSPAwQl/usHuGZTXg4ycUNKyCo24goLhNge2OneNy+LdnAOM0Po4
4QG//0o8QMvmvGrXWhoKZXPOsZbbFiGrUSY0M+0KT+DoEvqiDY5R7EG/2sFHRbHLiM+wdhfHuIKE
NZZr6bVa5PdDixoGrQnXm181PBWIsPepkC0bBDbMVN0ZQEGxkgsBGttrnjOEKdBtRRIoRgizH2d0
veYJHQw6o26SIR18DeJ3dt/rsRQVojICewb3QHLfYVEqVUxZ5/ysr0dao1u0tte30euJfgZt0qP7
s9OX64gR7+SiW+TYrzwLdJmMYVF2prPyXPqmJUbPucL++f1/6JP9q2ruhQPfd/WvO9evemxmmnJu
7iHSe44nr78HUd03Fws1l0wNIHZatqfHB2kMlJaYYzTLh3g9VE4MTyilmLC0kcFRpQ5p8++vfysX
agqFKoGhFeDVJESsZA85ytmVWDEFp40hqs48OCHHGaxcK01Bmt0uU1tuItAGlVtH4BjtHbKBBE84
iyms2WoPFtO/ngMsEP3iykTM+Ke/u/li2bOkBBA6tOmYR/zQ/nK5491mFXM9Oz106G3TJ7KAE73O
rFyDRjhTaVdJe7kE743J1IZ3pGmRfH3TdELKzyN+OlDma9dx5TEMpm6p0iz1GNblLUSREc5KZfb7
C6+4DAvUbmYctFtW4NjSpdJ89sFj0MTioQNhxhg3oMypFnVcDtvT/qS6TSWZq6p3r7uB6gcIltH2
ukqS0WWFHh4bvGTb2S7XeaDDix4yzqJwX0UuuZO1OSN5Xd7JaGj4/VgqjYX9eecNyqgs+u71P2/u
Uw25b/3VyzKi2UlpGC5W8wjOC+ZksmNXPNi7A20XxK/ZhrOodL5QpGH0D9KpFZhclau62mZLc9Le
xELxB3N9hkDS/Th4f1guqL1qS2pinJQPC/RzuqYJhgUrMoBW7HrDHUYUd8Wdv5ypRxPRjc28gxWe
FyOdlUgWCzLuPhY68sE0BdnJqPrKvX+bjkssXsde42+TzvhaEKgYdXZhPw0ncE8hILNT+yP8NTAv
kTOx/EuzcHr8XKd9jpqwLWdtXiasXrrj4Q2c47DfRXK0r7ho3ecNzmfGw5h1/ODG4gwqfmYQfJkR
OzvLyNBBV+pIGHO505N4Uc4iMrufc+3J4ki/R9/IGtHlKYpPIA7SRb95ibC46/ML5q8zz2wyocZ6
zPFjDwk6eWmH2lLG4mp9/MjfcpsY5ZCDnNSQMaeaMZfJnVRVriCIdpDGTfX04vXzVjGQ5s4bWQG9
eCzCydzToeEj5xiBG7J7GffSxSoDOK+/aetek6BuZwm7X4PUGZI/Kko1d635Y2weDshLgmHuAaCW
rg0hiYKdqs0gwFDUoNpcaaV+nE2SH3iQTLzNqpfFIMqFV9H6Kjpuq6+KH+3kqy4xkjkao0A+F9Qx
Qm1Yc9LWV15Swo4ZGZgJdxIHAb0hPLjcKQIoGbrPVKgD8xtohBKRp6iqFCVQIp3FCB8F4mTdj2+K
0KrPsOg0hyoS94uue+Iup4Y8rbKlvyHGCYRUZUAcLRTUTpBI3JljxFKQfXFxR2wlRzSGeWAksslp
zZx3jK1NatAipkwaUw69klvSNl6D1sdiA7tT+ye8bdDY/ITjJq8SDKe31U9wLVLrkZ7UWd9C3Mzj
ENi69Q3hueaqXvHi/5QfGlbsnhGcB4n6Qp+VzN8ve3WJKr5jEsgMNOuFeW2YreJtLOlGyHJhNTtU
xcqhNtVzBHJWp+iuTzCOIS1sUO8KgaP0MUtzCALYrNWM6DaLyi3+lJagdxPkA2GtOTPWoAPGaGqk
IKoGMYNhjc+eFNhJkNLPRcZ4EjOJjPGbDfUW1fUDix1Iijob8aSZBCBQTxjIwCvPQ+lK+CNGfxFU
LCOIKefYfFod6JRP1a2mc0ADy56R3BfVXuofX18Yl0HA4Rj+poFS9sfyq0rIcb1cF4odTuqzVK6g
VoPNb3QRQYSBVb6jSFBJi8i52wqskLKb+ehN9ToU30iT/dYbFwX9E18xwBJ0t8Y7jPq3syur+JW/
+aPwaykxEncZxpZj8hpg8pw9od6c3qflTDEB+bRsCWS+FqakbrOCRuhZyGvNDHsO9k/VK9V6PCQD
JfFRDicRl/7r/pN8KpqfYEuMrXJJuUxE93H4xI7GATAosnoGR/PQZ4MFOAzTlqyEsK4IvRa47Krl
vNSkG1A1j4HcVUz+B9J9DAuJIu8m+O9r+s5qCoA4lStW74XKf3gdhgU1pc2eOXozpqpVH/+sOC0A
mssjI2G+uwqPFW0Q77ekb8FYQBei/U1d4hFWr6QWe4AKL8blgFqAxHDSIPhVGLovUDhJtcmVwYrP
D6J3uQA95Rby7Ii6URjkBEAgK/RHObSnLfWISE3P22bssNMLLB9qmSdVKlqAq6T5bQIuZw2Rwcrp
O+tnsMk+FAEj9ZvAerWMIGbc0Tb9cKwnge+PqCNJ7QU8POW6jP36H3PrbCN+n/0p74y6PijBtQz/
Q2q1VflZky+vub4UpkFfiSRypfuKWwEJE41yE5/zFEdq9fq9Bvu+6QVKlg9Lyt+UlJbDD5K2lBkH
v4apML8r8q+PWRHdcFQP+OKjR1Hm2E4zEvoB+JKgYDEZzNnNZ7N4vrRcqdrFEUhM4riTIYfXNoM0
BEwahyMjZJJt02ca
`pragma protect end_protected
