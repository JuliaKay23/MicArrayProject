-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bZiRWg3QzvHLNW3/w7eaY/spk9jck3Risggh/ewSYwk+dGotHr5H8CeGgsPMakkZheggA8lCqIRQ
9PwSQ6/cBylJfopsXum37FyOms8qZRDti3px0GW8ncfZUQTnIiUpeTRJ2mZ8xivNCevMBkv3ts+G
KDgIGsPg+04PYRC4kSdtlgg22NSKcp2MyCvVkMRF+fFIv5SM6mX7q8JnIG2wOLjsn5pFZmqgiWSD
TuMPPWhJI/KBYwhOkqc36i+kUztkhvgRxip/hG6rTDEgd0rRBPB8C5zwYxGZsE/E/H0Vj9IwOP0h
D1i0rYwd84+gO5F45MRsUBtNgkCM8TtviROBTQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2640)
`protect data_block
PK7+ojYcbBcfUpwGiWC9+uuO/zWYoogWh9PJCrz8p6VVS9siPzHx8FtOfwKEv8uoWMUAcnInzUy2
GyAtralL+J2LGKQEEXig6Wdbmn/YUzccvTPb8vZu89PA7AdOka1scbDnFQIMWy8vmHrGMP49O24C
aUTTOqs6bB2hiJ+sNrHHC/kKSTfOjOrKYrrbD+GEdCYjbuIdq/3kIEh1WNawEA+wFaMOJiBfuGUS
wiVEnl1x4VPvug30WcGpk538caIgNalB1DQLxQwSodS6DnDaFKJVDRICsT3OTNQnKg3a4nFguMUE
kCpAd0UI+1i6XWQzK9et34qo57vBPrO8hqePvliM4bEf78KHga9MUKAEceDsD5VMWOJCPie5582p
MU4Y66EaCCONAlHYE3i5wQmMOnfSkUiJmOLndQUegpx50i2pHqGF80Ty1bdusV4QCaK4ZzYcsv//
DDak95iC3A9w9fllLVI4pPnFumc61jsbnI1RbjLZxu7SNQayRrNtGQj1lUZIsTn67sAyUUXOdx5n
/8SNuGteSrWaPCWufjMtqRF17vbwD7VoPhzSnglimkaQjuFi17nK7vYl1UhgdpApc6HD+deAJJcU
F2xAvXpyXK4VsDCAsVymkipiA7PibfSIipqGpNuwoIPwlvccSKkk22mCS+0hYLKJIUtMLQm3nqEh
oOhm9IEVFUToWT8cwoZEZREN8M7PigYdPTbKiWLAlqkgu1EJ7lChAcOvX528FB4hovREPA1vw0N2
JHJE5MCU7tvlZhpbyFUMHP2Et3Hk9T0dFwwmIMVKKhTO59/dy4CxW9BSjnKZEi1dpjNJivqCUjxZ
ryJz/hOi2pHnSED1J79YKXvgl+XzHDFHUSbFkeNC/Ob7+//U+cE7CNmwBC9ZTlniu5ImhvHPi61m
vjCA3N870X7bRMN4MsslyE58WGFXB22B78EqyxROlfnFAx5iQ0TwWGeEy3WYrD1wTf7K48j/OJ46
hgY9ZOv95D2zJXKTPxOKsZ6VtptWqgaquj727LphlAFFiOauKJRRffx6JBUhB7Xf+F2xHA+HO16T
6/LIdMLM/wqKfd+2wvtVe2Qgo6cBGjj6RrZA5WqPwPzsosrA5sgVSYl6S0AKotQcF4IwZrUt4u2T
SK6G7EvbOHGF+F5fH5lO6tjSrs4ohq0LjM2xIGLpUQbmbbo7R3Oa2N549J9ixsH3CiRn+Gdupki3
A/EqbKBL7fR0mLeBbQHA5TxZOqlUJ2I2WwdBngaakbGKtB74LiX296Ri4i+SRroW6bxR71Hvl9lD
qmjn/A15WZJaPrLyCURo8I24xxr+Thseexp2POb/YsFl3/ot/bB6pRSGQj/rMdFUnQXnJ3Q2TKAV
mWC7jYhTuAeDvNs5nFgf/fU24kQcvb8KDEDd0Fcnd7x80LNXQPS+LkqVO//BcNKZGlwyac3XrhtG
CCES6EsgbpFAktBRsQ0M+NzQWACj/PtRnESE3A4x5XjMz2pcIiYWEs8zwX1HyatGjSVhzA45nIim
9BqPqvw3khgFrVrY5BkmPIxOoli3sNKVvirbEgNel1W3km/PqHjewaexHpEofgdU6iHIgHo4pqNW
rB2lGUosS5CVaF0brrYTpExxqUoLq3H5Tky6t+siuwc2Re+1wGpu4q0i51LgcCmDvUmWmDW89aA8
Nfa+CoTZergMBtYIzqG7OvEWwVDg7pLc5jqSD2xruOQi8aveyirknhPNCyBng41x3OjcFBBUj1eP
Nh3Gyn9zvnvKjjuiU9ZvOAoqPzcj1fq10udMN6cqXHQZW5nzHQXfeL3HvuqQXE3Ad3N2HnXnA8Ml
mUSEjtAHFc5iH4HbOdjFQRX6mrWF1aQV+GSUNp+fsNVZIqhLRdKAcsqUF7bo9+9DjQ/AjoEskXGY
8J//IOYJT2LsklcrXydJpPJPsxmnk8ufDsWo2yBcBL5qJf29Z8mZV7vJweLIZK8sYWzwbY6O4TV6
LSAILQhjG0ni2uNqT3piQ1mg7WM1Xqp54UDz4u8IZceUGoNoC5WeaGIEZ8c8HioJm1i4SdhVVME1
3NznX+m+LZnJ+LMOFJcFNVZ0CoBrpscn/sDfsFTbYw80tvhYiFScuTBzVufHHIQY2jyWVDpLHuBe
7sRVbeyHyPuAVu8jSwUo2XTbndoAV75JgwBZbUwATdJJ5Rpfd+ejHvj3lI+07dW/bbSrRXbtnEJD
+kO/kHFmTViPvoBfPOyHR/8Pn4pONSvn3baQhrnLTos6Mf/0YyETO1VBcwQ9PkS8zjyQ5V7+2A0v
gG3oWUxwyTXCeaKigiPPG5tnKfRGVxyWHZkPNYLnO/kRpa/psi55UkxE6kA4GbN/5l93Kp04+xI8
nfTPfx/vMpUuYEOJcMuUaYnyTGz376ce4u8gar9HVmwfRUlTMzJVoLxxh8lsE54XSDbUt+Say0UR
leD+EXDJ+EK6Krz4JkHPgEvdi6Y0g8CgQxmlYR+J0KCXYP5zVCXfYAJfP+tM57LTpE8VMI/PiiST
MLWv+6OFwKQTH6Q5YNMHDVzySSp9OpzT7fNMly0fyO0k0NlrXKISqgQ6wqt/Y8NmgY9lQ5py+ceG
6oOwLJ2LOxa9fO0feqTlXjde7YE68Jza3Qs4aXwz9gxZgFxk2sgRATm3/yeR4qMmz0GgtXZicFIx
h+nFsVGUoTQyTehDYeGc7cwOLxYMkh2/gom9K/aWzr/WeOTj6kT9YWWNj9SNWwIEtAFNj+5HwYy3
9acwvJqewZBadQLj6iRo1UHYaAU2JD3dTLTwI3Oh3oL1m2RYsdcWTffNk3uoIiyqNuHZ+8MLvyZE
p0lHnw/uVbyU3l4tPB1CR8eRdcznHjXXer4CcECv+nPqU1MOMYe/lXtxrOQvBfaJmiobtjocFw29
n1RyFmUbH0IWcP9vKFNjvwhaBXZrbHEKLVhnCDVCYb+b6D0WniHIORSPrmqr89+wonLw1zD4AMKF
WnJVteAmhoPjBr6BaH+zygwjutc4fUnv8fBb03K8s7HeIWSmPU6/uNSz6uIoj2ojnbtI1Y/K8+61
9TOc0lGWqzXkjNlu2gvCf3LiA9c+JWbNq7YgkamnGaZ+1jrHpFYPmtLxZESmmzcytep5wI1HGK8L
k91XiEMWKfSkAx0XPye9satHGghl47cWyryzDEM949UvADtqAobuYq88RqNXy9wnEcO+KmM7AEn6
ZjvOXk5A9uvLGUjn4CX85xAZYvkoFx24CfXotfSiqZF9G28+ZJNsshZcS6rVXJa/26AM+X/62W3x
CtBrtR8Ao0LlHunioZHomB7mpc+z9ctFKgvWxD9y0EJvNrqHjeb99rZ1bIcotv8Kd0Pp6374uvbA
JnMSMcPCtYqQscSkcVrBMHJtp/Qw2HW3xKZsabF6IO6WSp+7dzAnLaMO7pXNXAm9ZDeSKpNK6k8N
S62wpqLNWHIXk4xKvxIZYFf5OjhitEtPCbcw9O5iR3nYZmAP8VNd4Q/oA73w6ncLVSUvW1wIcSfy
5c4b9L+gA6i+ZeacT/Rp18Zj
`protect end_protected
