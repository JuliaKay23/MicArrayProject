��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��y�i��6Nzywl�m}� u��Br`���k����O�{1M�1�*8����<�����Z���G���g���}$�)����$!��'�u�Ai����C ?%I=�Ҍ�n��"��;����-*�=�Hb�wa�v�8w��Sؚ-Գ"���z�ֲ��U������C�TW��~�揄GwT|]5jS�{��0���(1tz��J�܅��6��?5��yL$�`����5~l�	�
q�� e)Msb��(�}��T ��O��d�C�Ki�ѭ�o�])C:)���͡�k�n�R���G��
T|�U����e����i�p�f��~ز 7G�X!��@CĀS�$SN<��\���'r6�j��kY��d��&�����Ό�b�*�^�����.&��'�bʚ���b ���8��p���?��خd�+i\F��~�F�^��'r��"a�����LߍNHuZ�.�/��	8I��@Æ&�.��oܒ��w��M�O��V�J�{��n͋�z�i������\�ͬ[xB]׉&1�wgQ�O.1����M���=�,��D�޴ʂ�6��*�����M�)��3�o-�c#�O�e����2�'����ݽ���]�u{(��6�hst��vц�L�L��Cyf���^���EA�x(K��6����l�N����#���u�~�E`y��AAޑ͵Xp���K���r�o�_��>���kv(v��ܨ��'*��T�����n��}��r�`N������-��.�$�#�,����ڴ�s%�zQ0��}*"����@%1��EmK
��.2&	�{� �b�M�!��=Ӏ [K��ʴ����&B�@w;�����1��js��?޴�����CIͻ��.��G�而6_	���)t��Ex�c�~-fJ�@,��W����nSd�FG��f�>X�m�UG������q�!�EתF]�I0�X����vk�j������ʶte�<�����k��
(���Zc��Y��N�YT~�oy5B%���l{��)j&IY�$^,�O��uw��������dz"�	������.#�yq��@�e�W��TQ0�I�����X�j�t �.���-'E�� �f��>FǤ���T�6���G>�1ѱƆ�>�*�h�T���� ���������*u�[q�[�1�WD���S(F�Ak0�%�x�ǽz�V�e-M�^&A��ܭ��A�Z��q:�e�ǬԲI��J�8������-�&�4�H'�!��R��3� �D�1)�'ܯK�G�k��זΔ�E0��x�)w�"�LM��FSz������ٶ��|45�<�0U��~��B<pFj��~ҵ���>�R\�Xq�6��P�3�P�� ���ʨ���zf?�&��qAw|e/����m�Q�/%Ɓ�M�FB��[�3EO�SXTHl�-c$k���E� �D<t���8L��?7E\��W �ҭ�� ]d�w��!Ma̭ID|^5�o�KYS=n�>t��n$��oJ�Gl��9��]�{_�f�;'_��<�Qf{������.Gs��������SUs��oDS;�"��:�'p�*6�J� ��0���qRd���f���%�ɓ`ƙ��ּ�9��	H���]\��b�f�#��6?�����'��SOM\���Y���G�[��ؖ;Ix(���`�L�]�戀�M�_e&���\�<�]c�p�)�M��U����ձK�������U��$�����UD2��tw��܉�$1p��}�D��J��d�~l�B��f�	>�m|'<�K5S���l/�)
��g�&��4��=���!C�u S�dG?�%J�eC��ʅ��� 2#�]
�f�z��a��rb���n%�/l�)��B�������h�)���Ϫ�D�)�.�u�Ӝ�$!�yQ�bA�^�?���7^�X��o�	
3X��<�k������50�!��gop.�ob!�12�1-,h�p]�#�pN�ӈ���&��e@�s�=�˦S<��oHi�����d���������c(�1r�2��yl��n
Ī���)/��\l�k9�9�J�!ׇ�<O���Cp�
&�s6t��E�Ȥ�K�Y�I�m/��>Q���`�$�Y��:���)�i�9�{��A�'vhB�~��"t�ږ�a$���3.��k�[!�ނ7i��Y���{�v�r�o;�6�Ϲ����"�l�?����e���;/OT[��8�[�
ӠƦ�	^[�_�`
�
,�/�0O�-�c�a� ����O�P��I�#Z�8�X�ˏ�-�ބ�`we�IV�]��[���\�.����,�(����3�.�1z�B�`�,ŷ�}h���xDR����h!���ڗ��!�|���7��������ʲ(�l<����a*ܑ��}���;ӈUN���k�'.�N9���\FG���O���4�[� bJ����SL�4��Oݛ�l5ٲ��j�yXN+��&)����me�E������EC{�+�|����^��Y7Ln����1��c��7��L����\�F>��$����(ќ�\PB�Z�B�sA>�ϲ��(�ۋ����I��*���^���O���<�e2z��b��M�(��*��[�k�9�FI��X/�I
��j��Y�DS7;&�������3�o��L��y���*����_Q��l+r�8O���0���m~3T��6K��4�2�A���H�_Xf��J�U�7q�3�ا��V^�,_�Μ�`���77js�WmY/M��gG?��y����>��J��'��Y��|Z�t�UůS4�T���ñ殯�_��_R�f�6п���3�d�R�ꆏ:nm,`���Ht��)�]k�T6�N��U����i�2�"[Ջ�GWv5�5%�S� �W@k��U>�`
$\ց�_>-<,����<F\�:��4��?���>����p⪫`i�W/�/�A��1"V�M�m�M��B�	pŜ
����7�~0�9��a*�mE'��7X�C��˜�����R�"�N���1en�j��ri
o�0�`ǖ@2��2iBrs�`����K8J���e�*�5��O�E����m�A�7"�YY�BN��m|ywg�Њ^<ԧ���$1?�"b;�V3p Խ�6�mf�b�n�����]����$<���P=���+�4�B�D�9���*�<_!Dɾ��Y�=�����ʱ���Z���^�~�j2�\��&�u�
��sx��8z���Ǽ�q7t��:��ς��X�[�����c�yg���F��Q���@����救^=�[�� #B�V;�?G[�Z�������3 ������t���Gg��3���3ؘ�mI���T�复]���޺i�>�i���lvy��B�2�i��sG��<^�<ւh��߰�~^t W�x��3r�VT��Yʨ����w]��W����𚼓d�<;�^n�9����M��-������Q(�޹��������g7�;;��WG�e<�Q(sn�Nϴ�,98��U����*�c��Z(I�d�{����k�hA�cͪ��Ȭ�J0�W�\����.��g���Ø-��+#�"�[Vi��'�HB��k����j~͜`o)��F��̏BR*O��Ɇ3�|�)ꞐϝiRc%K\+�rze3��3H���v��Q�hU#/����2)j(����� ����X�"CDY��� �O�W�#��sS8ƌ/���3���D- s�����JG�'�5o�$��<��.�6%/�vC�J<$�`&�����k�0`=G>��`��	i'�7��m�yӒ���s�jVX$�[6+K=�$�ѧM�v	9y���>Hj.5�s�����d<�:�2�'� {�a�̓q�u^��n����̐n�+���o
F���"���:3�zq���yx�mL���1�.�WaȁLy�=3.U��=l�I��)�B���S��;��NBl�j�k����uzx���4B�1� �;n^��	�&yd2��D����6Qք���+d{ ���8,J�	-O�(�5�C+��?s��!Ű�d�r�.\WZ���&�W���gG��'60F�Et�v� �!��{n3��,���p�	V�M�SWg�1%i�s�B�ܧJ�vL���8M�ϗ
,������x�M�}j]8�A��T|"ѣžg��,���Z���!���T�ybg�,�-�N,���`���	u����;Y���Q*�u}��ZS~+t��J���-��`��.u!y�K�Ý?.	g��5�+T�4����d��	�Ռ�����1��*1�� �ʸ�ܪK���n2z�<ʎJFu}]�OW��8<��fSum<��|5p�2b1�1 �nH����v���X�L�mdt��mC�?!�lKŋIu��Y}1@1\B�v@���:]z56P�������
�c�T�N2ߠ��Y��O��1��[�z�&5�0��u����+���qp�&p2����o��p�����G�
e�5�X��Q7>�E�q��SH�
ٮ���"�H����(�d�����)!,LJ�W��2	]6xCR?��w�����M_��w�X����8��|�QL����z�z�޸���?%Gͻ5�<������Bj��0��]�V�<g��w�4)ė�~��l�A�	�x���m�j����I[�_��md��r��iLs�{��8d.���o���ܙ�Q>��=a�W?i����j��v a��|��ޟ�K�7�§��ۥ�~��0�Ý����s�+�{��w�~|�P�3��	�<25L���yw�K/�������c�'~\�����6�I9@���,�d���d.�;�z����+�� ����d�����#I�@NB�>G1�7WJ{ϓӪ�r�a�B�pʫ4��D�4��җ�I�4LINKX%vv{�h7�c���}��Q��}���eq�'�
���BZ�� �R�r���6h��Xߐ�|���Q�Lh(v������WMb���@�z�z��5 �_k�艑>wr�y��y/K??��D�]-�vJִ�5�*�c=��h+5l��Zۙ�*s��0��ߖ ���G�3L�m�쿭���1(�;Q
2��jM���<+�V���)w�ݺ�9����;�I��7�`�w��q:7��w@>�$��Q:�N>^�]U��<S%���oL�_!`�0⦽z��oF�w(r�X�H��4�[�2t�_z����%�4�4O�D�~�Z䤉��s��B�������Rk�~%)�Fg>{M�d��!��Б�D�}GT�����sNE�g9���F��Oe,"UoDVp��W�Y�����Da� lc�����rUT)���.!�v�|؞��vBo�|Q��m�=�o1�A&�zRq\�Ң�k����J5������s>�H��oO�#xA%Ŋ4�g�p�q��`���d�>g�J� |mpH����m�N�r��l�"��-�ݘ���Lh`t���1����q�,-|��d��Pȹ���]�y��B��/d44"Ŋ%'ͪ�kY�ƿ���3��
 �x;�,�aYaR�E����zF���G�C�%>|LoU+qv���Q��q�:�"�G$��e�����4,Ks�?�ދ���.8��\K��q_��-����" ��*lÿ�o��{����'��^vn�^+�smmj��ະ7���ۍ/=N���rL$f�����֞a�: f��Ϫ]��4��F�������D�#䑃O�3��-��Q�uC���e�~��+Qk��v��ł�]�G$ŵ�2��[����K2˓vĝ�Vx����ۍ��·��"�C�9`N�m~��
�絈�V�?�h��e��U�9[���bp����~����,������z��T<��4���,TWS����G�̽�?�*��=�Wb�C~3~Q5�z
�~޲\������{4B�.�� �P��H��r�V�N-,�������r^8�vL��s�����%L�f���>@�X��oʰ��$~AH�ku���]KӍŀ/���L8�G�*�f�Jn�w=Ƃڭ��U7 
�k}M�_6q��������i��*,E�JI�u/�.�)ۗ68w;�8�&w��|v+�N���Ps�w�7���U���wJ�*s�NB� f�dຯg�!����E\�kl����$�p��aw�y�E��Ը�e4����Y��1?��e1hd���r�Mm*,y,���Xw�&�����R�s�$w���IG��U��F�������D�q	�W�?о^�MEɊ��,��z��
�Q�\��wFi��
��e�_��i+.5����%��+�;�a%Pv_0,~�L:�`C��ss���Tp��