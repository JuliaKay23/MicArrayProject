-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hTtz7mXcTMgOPcqcFJ5KPPoOsSfnuVuxYHY4EWDxXBT+NEel3capip9TL36C3IPqrvWmgTskc0KH
rT667k9EJEvL4zYpaCAlBlGLS7Yy6z4usIsp7eNsvcYJmIBLJesHOQc/VqR8RMUoB4dIOikJSQvV
O+LWJQj92izu1Z4lAQEQwmOumHmYKj+yPKwp1EaAk68hL/cxsXawwlobtZ93O0YreMhIoV1lGF60
CBwzxapS83C5UbD0G2eFYbl4td3iuPHBH04GjrIGh8ChmG8n2qJyz2S3Q7GuPfSuZEeMXo6NVRpv
FM3oJsShmmHdpweq1Ub0ZYYNPtaKB9YD+MWLNA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5328)
`protect data_block
j6FFJVbp0B8XZYi2pUIbZheG3PUieuriE5MRnEjUYTueTBp+mBSnhkQ6OUFeTs2jDBKbyDGlR7x/
5MwdF2qst7EDqd5nt95kpu1Ov5Sy7/Oe7wxKf76o2/hTxFCF+FI/kGpZPo2nVE/D9wPzmKngKOV4
UVsNlr9pIraB2xrV9CC0rf6cGT8+E75EQckN4l5oDHutmvz/k6F4CIUDtPnrEAEgjUd22engScH3
gl5sgdN0rr+ReyFnDJoQDQlVXdAiPvcPGllqeR8yauHDHcNYVQjJkV0DPbNDM9+YE/RcS6fBrecR
9ZtSFgkjw25rQs/4Wdvs3rjQi1XuxFFwklu3b2tw47mLlAcRUBGsqojamv275AOgfJ82v/xNIfy6
0wrLB7q5gb0DIZsUFkCfo3bkVgtp0GX1M/Tc+aZLdq5GGBz0rwY2mTNAdvefsLgB3dpeIoTXwJjU
0dZwi4eqPWkEsygGPqLF6Cq01mp2HZsSbcdgWCG/HKl7TQcFvLUaBiymWrTNycg4GfawtG6T2Ef8
CnsKeYTgHjg3AKSufnufJAnGKDftydwFg1LNi/j0KlHArklayHJkC75Pu/PFBqvm6RzLHDkfwYgr
PV+HcSgZJ91ZpOlIHcOeqvg/A36NG5Z+c9izgNQPhwGg1UgPsAr1D5UmL60E7WiMZAuc0x02GYQc
hJH/e+lUAw165l18iV2gBY4LoBogRNZxNQkRKexADuv3cY8fiEz8Yp+/IIUOiVs2GyXERuSukCWo
UX4Z3+EOsEJIDJuszMEAw8l6LOULqcm0UBws1MymN5+wX5HhQr/c85W6p7ZlsJ1VnW2QlgEQrcC0
WcR2/RA4PqHp6YH+YJgLEDNV0XT4KCmDVdvERnICoz77AAFh9M5ux/+bIJnkzetH8TA4pK+jeJlO
X9MZf4Yom+l9I2tdsCLirQ7o4Jgeov+UAMGXAKz2Ud0Di+dXAcUwrBl9IlI45h2l1RIQfEdnnbEp
pbZQH7lGQoh/MuT2tIWc1suqr5xzvqAoO6Z1xse4Qr0EhctlkSzHs5vSjsQEnzvFXJqLWVUEfDtZ
u11tYQHNHuTliqvyQONBh0Csf40RqweN99YNoXJAmb6x79sx6l7P4lPEu4IzZz18gRjeR/aU8JVE
ji18cwA8mWQVOXJ5RrTVATZS4lsfraUtNscDqTvVPGIjx2JMIXqYGeGQULQD3hIpcjiW6sFaMNA4
uyZkIjF9V9YoNOuim14R2mUWQ6jJDY65JYbcK3Cgf5U70q5N7/XgF9/XCBrTz7bG7KdGXcq/RHNx
RpNK/N/s9PcQM7BZIhY9c3OdqGS41YY+OENnIfBkk5Z4QAyNmWLZZw9lQ+OtqJzDXzcVkbojsMgk
+i6dhyWIXfaG2Aaph2l03KswpmKtwZnip80cU28ueegumdlYwG/zEV7xHHiC9yTToDdkpU6gy3q5
TDehcpYMQuL2bg4hN5rxIMWOvy2+IN64KPnAn5fvzfi5EjwYKu8oMl0UFe3OWWHYi3N9cwJRN3QL
t2eCyUFsrfMeAadeOrAz+FJKOW8gV4Fw9pGoXIk56O1s6c2CkDyCkSdHqNw7DXWpxvAYNh+yaMdK
E+ekFgNBddsnjFAQ/1HdjLcqbrNVW4fS7MkYTNs6LQhpLNSkXto8tXAoveELu/R4Dzt2wG1HW+nx
K8Foli3nFnZGMWY792fFjcUNEJZWc66YIP3sfNqXRFl8RqSpxnys0zri/Uk2X9LFLjB+iLRJ41lQ
FjGSZNp9L2LPyM/RvrzAN+amPDH4Oz7+RuxE0Somi2KXH1VTKEb7MRdG7fG0vhppdk/t4yOxbZ7n
fPOnYMnzyVz4IhfdVs1QYWC6ma+yEJHLRxkul8+JLrJRNop7N9KIGfpWID7azCawszE7VdI7P5+1
3udPVci32WyZWYW+UWt5cv6Th+B0piNH5G52GE2gq4OpnNnG+63ifWlArmEchz4IbVbUxJu7IKtC
jcemTJ2vd5rHKWzvy6CZloReSgp+qYBf9Y8RgAd0KOdAqLv7YW/GK8Uq11y1+kUud+SyJ8QnlTmq
42Df0v+8XgoGswy75lWQ0roQaED4NGUsfb/IJl/OOINubTdI3zPbY2xBic0g2jsjsXusBMOMHl+h
LMa36/k9reAp2uuqNAwMGhP1o667FyY/1j1wnxEWTZxeavRzOTf6QRd93lelFsyRSJKOryA8Ph/U
V+1zlxkE3CLr767Y02/qsbsSQ4AeKrtLdRXrIs/V8J2g69ha4ao7fR4bqWJYmByoQDfLGzI/LW4L
kC25uakFe+e69cCAleQjUidYjHpVqFzXv1AOuE7f2jYSIdajODqFV4pQaFOADREQaFRpRiF6nfyb
UE275/GGWev/EE+esX+qTb9I4MLYCcECvAX3/NU1EQxlQWcF8Y+ZVGSr9q11oVi4n9I9n3Sg+woD
cxk0xHrcF4yN7tuxvhPf1pKdf/sLP785hkLrWS4fFl1iJ2Gs5tjE/Pk7u9NYr4JhBgWSytUv014L
N/WGvre77fGpdfgwp/557GBC2yZiUiLkWqDOFUogfEwoMvCBtw4s4bCTRf1PoSMFH1wZ+j1ngWDy
Bsm7b59Hw34PcxECCZUCc7dxZShEtUliy++rj66cCi5iRJLE/6ZvzK5HQYX/SFIpv380VK+encqB
j9lX7QzxMH805XHTaKu9YplUHCXYZRuBhggHSMGboxl6s0BnmGoMG39JmmjNxQ2ckHBpNoal8N+h
wD5FvUAHDEEiEaw6T8TW7ZlA8ADOdlcohACpO4Z9sxOX6oPg276BHFRk+03zHQYzij0Hwm0GjN5N
4f9fR66PsDt5yBOXIANmeoc9+Y63ZYrHFyuksrsOme6OFFkYu00ijvClbVc/DaCD8bBQ2oYr+S/V
iuD8B0Zz5i5fFclOrow0xrIIMg7mDzeBvGdjNABFbPPRKbMktB/pnhUM9HgEV+rQqRMhrIYUgTTs
uTHKL8ebpyxCNrJ65pwDN6tGt0ckS1ZTH9EoMVy6zsazEMK86O4M7tslQ7MsP8DNQlXe9yCt39EP
EMArkv7GKkigJXbGbutLePgkNrJygMW19+kB1zcWK/3t1NUan17TSUDaZoepLOZD477dj0YQ9X5I
IZWJF0osuQ8/rGrv+6uEuQzTXlAqLfmIQyTTcwo3yKR16979NG3qiG02r592cF+MHQ8H/ML9FaUg
48tK2077033JPN6hfGZNW0zPO0mybMimWszNivBZoZEW3fMJBcsDnImVSythv4jaBGsHyXcZa9Wk
3UCt0sOitAAevVuAUfDlgX/EUyvH6wHOevIStGkp87E+Yc+pAkyz4IfNSjRw3tm9gO+j21eajF+y
9o0gmUgbOPj6BtsKQ3zjqtviZMyIhYQNQjyxYPk/2t4XYM9X4vqvtl52xgJRYdjvX5dBx9VDOA19
R/bYP6YXaV0fuv1nCALG0hLzfsRAtZ/im6YItqmAXnt80N0YNf8aqkamPpvoMqROlzWLnCSrAuYZ
NEPt8hZJhw7dXZ4fhVQ9yGEidU6YUhHqg/Q+vZ9vwCE8OVAsmhASVTE7ci33wyhN3wJuJZQ/cL/r
6aQrhozsXr3e3PXERLajSce6pJkdnVg4ml2vsXmKXvwT6t3IvDHy0Um/2koTHqDOcLTaFwzfE+qo
sYC5Lv0pA5Rz8fr63QzCfofWViiWhK/IAFj16HI2qAH4wlmizZiUvLdl9ZMXMuYZajhN7xpejQ6A
D2SJBHWOhBzxQC3LxtMJanvo6fMyYmjCtRRW8dVLPF++RyRZw45O9X6X11HZQswhIuULi0vRAR4K
4qHANi8wKk5IPWuZOPD+zUwtMBWq7CoPKeNhqE/Z9Z0Ys8d35fTliyYwPuSee6mePGQ/JD9xAC2Q
+FeNr7vrGTdHLVzIV+i8jw5Bh/JKWiRKaTzu178KqEFQ/ZZiqGcmiBJ9ZATmoZ5+DytdmgakLSyZ
yfrShPBvW9ZoQPhWHgu0iC49toUfExC10CQBEZfh7U/nK9rCdqQfh468lkb0GEC4YZxeI2ntZXPw
IMRWI5Atp45QpZlxh2d70eutxzywWzAQkCDBdlhI9n5e9cEEQKvet1wLv/MwMan7EqybKFp9GXex
gWcgtgyjGBRShhbMqB+mpRSAsj/NnC6CWnKKxwPncU/kZTH7IHKmtVfd1PHPVpVbrsAxVxh737F0
4dMqkRkxV9+vy0arh4P8XpVxafq+stBAZW9C85Ztb4uT7J0PrREj9agq22YqOrtPvapUkMGC/BkG
lQ11J0ksGGDE6Q2ffFI/bHlgCX8j3ft7PjCBWfI1XEBftFXH6VgzVMIE/u59V/M8BWUnpHtB9uZu
LGEhpsNMAHVOZIlkIR3Q4uyWJ3tyFSmLNG/9HdHmvOvyXPUxGQp3eMDfNyusL3VgBE48qXYAHTfF
pCGjmAUfPL6XIHWBvyyszSBVor98Huj4wA07TOjtuSmkqFQy7AOagaAMB6nSwXUY+h2e0qYvxP/L
s21cLHBfhriXyBHyLmF60gnxD/b5hM/WnRR9t9zdAK/LYr3q+c+9bzIrf/NmaYsnVbDJQeHdFm0W
jzt5yC5+vpGzR9yduBWvER0v/+I3GXBV83TBmcdMldkDQ0bgacgEn4luDXXL3+O43ox3EcpA80LV
w++xd7Dt2APs5/Yw4yM7FybXTjM6mTUyCkZbcSRwnPGdYu8zhkyzsBjEvjGxF0HcW4INDpdx/R/z
U7CHp3gCkXbLGDMHabTwnKB1JNrFt6ckGGkwpQilbdpQD/6Co+8Co0L9hNyKLZr2WMQdWqImHt0p
MfSybtC2wCqgBI4Cfz+zwJNnIa5miANSFSh6FZdWwNVqC7ydmT+8ftkbildRm93875sKjGtx5JUX
B7hXa4LOUqpbkx/JEweerfoZWD26j5W34v9mQ4ynqUSFUUgDaRbMxc9tdgn63l5PKSQSuhWEqKWD
A5k0nuKvEcTdYkOi/C7JdO0w0o4u6LvNxrh8YCHDmu8pEFzlBCvpVJU85nD0P3lG10ls1mcsSnsX
QiiKysVUxcAQNBoUPMY0928G3RLqzpJROyTuMHl+/xydXq0Mx5ChBfm1AvEiN1DELQ22o5Z8iomx
VWiiS6uXlONAP/vsPmvBxzoRupGVHb9oQnMeGWoJBJRBmbbxFmlSp9cme5gPi+c+Kf6jtHMvjcv8
bX71LrB2Z0R1sGQ5CAm0NXaT/4QifGSshzWAEu86wqVLrSrGA+lJvIKxFA7mif+4ws/qEOZ5xyuH
elgBlraZ9wAkJyQgRk6lkpstp8aHH2upGHeXh7y1ZQ+IsAD8vCNyj6IQwhv/FB1V3V8A8QfaMrI6
S1xDS/uwiUQaWwxTlrRkpG5YQUMUu8mLLfK1FS6embIyGztHVPD6n1Yd4ZJNZVHGgxdIIRFXjt2E
Ke6dWvRL0QNpATTYSiRO1uRo1/ulZuZPpythsZvZlATVhF+dEBx7pi+kBeel+AOji3q5Sb1WWr/V
jwMdeOSh1llF5gzSPnThxApHsE60vzrQcJvEvmpm1oqgZqd1ouPkWfvTZQVTyrkGvPDpYK2Ae2ce
0sHDxP/UDkAQML5k3E3ZLoFmEO4XWAmXR3+yVJ2mB1bljioWMX+lBvaObHCepWg0oMtE5MxA3wJy
SsvMSL9hsY6O//gw3fZIf9VHL9rkHMja8ZhqvKXwE6emwiz1yOizeJ2v6c1I4iiEt8e36qeookmt
9XumPGLj451U1+WkmRR13Fv1tUBXbuvDGZhJ1MwzCmsJdqxzo/PC/FnQ2wxP7pnQrXP/yE+2pSQC
/0dgH4OsEqu9k6gWW6tGCgS1FYSb+iWUbMDoW3AOpxYqNGuHF2l73r5hqu75Z61QSA3tL858lUJi
8DMnhM8xNUu47mL5W+LCrHBdMwLELeFSOdxTidl6L48CYaZO06FZXDP5GCySaSjssrCAqiXZ1wLv
x48j9etpqA04JJ0pr84rbTZV+SXN1gWwrxGNXGXdSGxycz3w7SINKe5r3BPdk70y3L/OdAuANqbv
uC7qwff4b5u4hTwgK8+aBe9Xj4raPiLDi0Zbg+bz2chbpAtTTFGv57i1Pzz1dkPZMOBV6LFcUbQe
dsmOdpyNuosmGG6i5CsqKzEpxQ/26DyRECBxdpv+SGG2hF5ZyEZbUghpysDQHXDSea14z2Eo7mlv
rEtzjkIf2YqeLsjttho6EaBlGEQuDwaEdewYL6gg9MZjIcZEGMpQ20LWqXyPZEQNIKBUtEQLlnbl
oLPqg2ismrHLTePcM0UIfB64zf6z1qTlpOGjeUD6B0yl2VzLsuL4l5zkOlbT05Jk8P5aYUXUnzdw
u+J552Tinw+oxkHugvoWX0f3ECTeH7kjghyPE79fiM0ZILl4yxEQ7RipmFS1fNwSpPoOEOvtejM6
yt0GtOvd+78c0Kir9VUqD4q0okPPGItWfAky5NwhHQTlPh3ngMDWdPuoM9pFEBIpRdda91b2qMXZ
wakg1IPM6DWbPQUkkq+l5hDNs2qhGWlVp1xhZy4DisFsfpVKERlXmv2IHGXUx4jCXVsw/VZtkFjG
d3DCdcDJeygvTeZRiAgNP64fTzuc5OxGgkTYs94Tsy1GxmBLqaPC36Fc7ZQ2r1gp8oicb9ba9Hvi
TWju2/si9wPep/748wQxbZHmYKnESA9CjwtUs9CLu+sVur+SuOXK1IgdjUDoALDu2JVmtBP8g7tt
Pf73QQLJWmNVFbNTKYOv4q46aBoHS7rEDTtjeJch/emrQkfDC8v4jLmhEYVfT4alVi90mpFTMNff
otRdDoM4cglW+Sa5vEn+VzaF+C/c9rqmgNmfG/B1tgRBUMT4IMhbCE6kNFdPxP7jLc/W5rsdlDGT
SsjRVubpn6XoA/SZhQ1+sRQgE8DXlX6ZQaLMJHAI2NkAJLQ6c6dx3b4J0fZucpropnPjSud0vw+5
3AP5sVwH+WccsXw19RVBReu5RCBR8QkuVZrnmG+bPuGyNfoHrfkgksEfaFaiwSWPdBVO6dYxwbRN
dcZmwA4nue4etwGYvxMXx9AhJPsDeovfAyEmzpGs8cQ5YFcdTdZz3XuFsHsuMZWAkqYpv9Lq19LR
9iT5dJVb8o+lgG1AmSYw4XbaqBT0hjDitP+J
`protect end_protected
