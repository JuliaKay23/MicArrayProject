��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�GN�Џ	�Uy䚜cs��:�47w�D��M��b�����{ad�H�Dk�ªJ��^�|5�x�vy��B����a]gQ���!�K�u�xt�e��4��{¢�H1c'��TsJB%�Mt��Rh98C"���KFGO�����So-&��wgL�v��b������I�6w�p,Q4��:]��rptc�0Vd�gWw��*���T_���v��S�>�@�}�)����6�};�ؼ9?}�`x��T<�M�(�lv�/1;�X[eM���'g�~��n����a>C��<�s]�J���i���H��I9�(]A�8x��H�4v��t�:�%�臔+P�[��t�����yx������L���g�Z ��4���hng�1{R%k����c�~�lA-��d�7�v�~s"��)v	��%�H�|��+�n�d��cܜ�O����؅q+I*0���6�����y�TyU���k6���,;	(fΪh\����1�֨����]y�,�n�Ds�l�l��Tb������j����3�=+d�R���B��+s>��J�.&�Lj�q�kј���[y����,~|���,�=*��ba!Iv�5�BȲ���j%�'����=t%��l�nZ�r�}�&��	���֜{�T�Ը�� �TS��A>xB9�I�K	c�����L�wk�����W,G�us��+�+P)@):��s�%-�C�/����V��6�0݋aQ�^'H�	~�R�-YQ7��\}�����I7o���3@�΋o[�����j�$R��i�v|
�Ǚw�9O����S�%��yh�B��.���D��B6m^��j{���M輸y���%�x��Ӟ��QW�iH��7�UXx�2��с�@=�;/���}�~�����S��_'G����
|�πo(^�=UyQB�D��\J�.U�]
�T�>vF�Yl�Y��T)T�DF�����.���B������d�U�C!�aW��{ߊL��,�9V!M�|TO�Ӌ�<Z�����?��.�c���4�� ����rr�8*0@�{����P�嬃�>�N5-�(������Tf�"��m!�@�OsE���}1im��#/Y�h&��Y9�3%�q;	��@���3�h�ĂXj�S��eE>��װXh�H�(�%�	�&��p�|y�hꕨa�J���|l��~�u3���I-�S�b���s�O��1�~2`C�5���^i�!�����P�K���l��|x+w[v)ê�U�*ѳs��������5�<02��\��<u*xu���!�!�1ˊ��*g)�}sR�����%ǪșΏ�H�UH�|^N���96�=����T�f�YI\��=�����k���� M��>x=��gQC(κ�k�l@\��T%湉�2$��ƑV|6����%c,^� ~�x�aɎQ�W��C�0�*k]$},�J�R���̒4E����b�@�|���sr7Ԉ-
^� ��m&��A}<@�gͰ����4o���2yM�H51�2v����Y;:!�^�q�0����7x��e��cl�`��O�bJp6ԢD"+�c_��>?7r�͋���1��׮���"='�y0�f^�y�Ft����9C�_����@�i��a<�tTR����,��X��.�����Tt���i���A��.���tߩ_��VC;��������h镪�>K/䀹P�TeX,@�Mq[��?��w���'7�@g���j$Ҋ�y���bFy�մ`N��������k��zI�Ga���
hIܴ�4Բ���LUR�&53c�K�A|�ᄯ�FK�xr��%�(��FL�g�M��u^T�����:��P߯�s�7��]lWC_Q4͔J��s!�S�����÷&�5�J.0}�fh��ˍឤG��a*�gR�w~���z��?p@5�y^ä��r��F�	�z��5��?)aqk���݇�	*'Rc!_2�q�&���ߎq|n�P0����#�B��䯂��
�6�rU���-%e_]�z���W�9tCd���	q��c���c-Y>�ŰBt1~V��Q�P�#��;�:�H�!�$@�e'wʑճV�����T��N�kU����`I~÷��Xr���m�c�ڟ �k�wIT�>XQ�+�}�(t\3�<�ɽ��������,���EH�)
(>���IB ��}��h�5�>����WT�""�����=���5���wn4��Mj�!و�o�"j�~��8��Z�|��w?7ŷ����~���t�{�	�P���p����y�u��9�����9�ĚG��&��K�/�k�]�(�7��w[������sQx�9�;uI�?�Ӵ�9�������tãJ���a�S�0ݽk�[�� �PS�YC�׃`�5���v*>�n�e}i��Sm/S������B��y3w���u�B���Gç�%��FT�g��JU�^���g$��W*u��7�G����4��(I\�V�C�8������3�~0.�E/�n���*m�.���)/;鋫��6Ro�H���4���?�m�=&��!9��/k�ې"�!�L��NO�G�W���+]�hN���yM��+��D�����8���nWz+����|r�ۥ۫~�Po��l���F~�#�ڔ_If��������g��P�Κ;�:O�f�����EHn�TB��]��T:�<nJQ/"$Z�Ze��?�oX�s��+�S�m�ß�����������|N�㮡�~u���'i���UW�yn�6
'��Ν����t+�`�]*�@j9�����3>�]����x�|�����n�>��
O�5�
4���Nd�!Һ��Γ[!M���:9�o h�5�}��6u�W�y��'��e��ʋc~�)���-ə��k89�G`5M�(o���Br�SMNfx4����gI$���-:�~�ICd���	{�(i2%�`���Qy�FQV�B�y*�)J���a�EL�C���2_1LM��'DNB�Uk�X�ȝ��/�dmTP��%:���=�P����B�Z໪Җ���ѓ�
����F~͠��9������H//��D�&|F#m�����bj��$^w{��Vnxs�m�	�����.�kT�f{#�=�4��0<��@�S��@��of�cVvw�Jn���;#�@��H,�p_>m`r���	g�S�v�����h�V}Pf�����^6�r��An�eS��g2y��|m�l�X�_���<�-������
u�Wˏ��Ҩ����E�gZ��3��}�a�p��H*�P5�m(ؼ������"�>y���)ɫ��+J=6o�m����߬�\Ůr+m�������&��;Z��y�Γ�˶�RV������u�Z)�YM�dJ�GH���F��M��?.����Pdf=�QKE��Y�П�=�&e\<Te�GB�(�K&\<W:��3��v�I2e�@j�v���i��r���mq P��W��|��p�\�c�泈�������V�|���k{��\�������Z���¦�;�u�6îs+;o.(=�GH�J��Y[-���ж1�E�WWWi�Ȓ�w(�8/�'����8��ۋ�\��o�aE�=�������"��W�ǵ��,@@�9M�*7�6k�1����\�Lj�-TˀT����g@*U촨��Ш.�]�?0� n�L����'�>O���H2@��1�Aű��ܴ7��2�t�Y�9�8w?�Nu��I0M^F�CĠ?��d3Tࡏ(�� [����"^QNs	N���G$k8�,@�ۗ�Ѹ"�S)׽ˁ�8�м�D�#2��xT�ݪ�N7jL���E���z{c����8�A�����};,b�bG|��i0��	�����[nU�}��}��e�:�@M����9�Sr9\5)S������e����>-����/����Z�f����rƓ�k��vKUAA{D��#��ʤqPq�3?�g�R)-"�jHxK���p�zQ��
���M����@�s������g}|�����\F�I��Kz	$�'Oꋂ%vg[�n	��l���v��54��N�/q�;s�_ar�������'��f#^(���.-d7q5�o�i���=��)a���7�;o�0�0z9Mg���wNn~���a��]��:�1��~�S�-��h�V�� ����s�q���-Vq�5��sͣ����� -�1y���F��ŉ_$�4!�|.��`5+T�z4����<V����oQ]��b�!Wk�r����ֿ�=ߖܠ\���e��q >�4���;����~z�=e�s��x���^��pT_ȝ���s��Gs�;�~�<K~5�+-U�ʬϹ<|��N��?�l��w�s=*�u�J��s�>��m�ZN���?*f�CVCX�ȻG�����Cŉ����ao�<�E)z�����0)C^��,���K(B�E�5���6]���� ��dq�)xs��'����FY0��JX%}Y�m��%�������#�k��jI���|��@�0l G5ǯU��@�%���}Z��R��f*n��B�V"ظ>��k,Ӝ�A��-Y���t�����cw���l�nU�7-�#�(��b?��XJ(/S ��w��M�EMu�8m2��g?����*~�q��%S+f;uA+)ˌh��������e~c˘#�d�������>����*��C��J��6��T�J��˔�M��� к�R�:5+m���(�qyr}�	����8������������jC��,e�'�Zx�������8��>A�Y*�)���t��Ys�����K��@$��\ �c�G��\M�4�Z����e�k�'H!!&1c$�,@�$�������Y����l4�!���[��n�����������&��@"��v�!�f���<E>���Z���i�SM�$(U�=/V�~���8ͩ�S����mNu�(׏�XW�)�7�>���F�A�49������0pMF¯�O���,�ĝ�F��~~�����Qp��@K��~ߖ��p�Tt5���l���FH;%�UE�\*��u��i;.Ӹ+I�ߘ���R��J��v��*u�F��N��T͂2���:ԙ$�r�7�"8|���yuY���b���^:G��mKS{�͓���ճ~��nm_����DD3�̵�Q#�����ʝ������V���bq�o�L������!d���g+�U���:�K�%)�֭���~��!�Њ�����b�3�>kv�G���\� 얽9!_wR0č�����L����*�'Z@��I�)��� ��q�Ûo#�p�y��V^��o��P�^<�h/����`���(��W�T7���l��. ��VEd`�y��{�)�pƙ���I���y��>��$b��[�'":�>XΑ�V�	˩M
�@�ު�1��<�o8B�{�8E��46@.���*{�XY�bL��Hn�T��O�Ç��!804�{Y̶W�N��3�8����O�&���*�Ns�%��,��]~���ц�xxN9�1#���A�	�w�u��r�F��#y�$7��P�*g����Y�_�	9�#Dˑ�+Q�mg
qm(�%;b� ��d������}�;��v�wl�LL�q�򼇐 ˕ �|Y9g(�F=x^�Kd��w�|V#��L��5oI2A�+������|�4���j̓ϹH��k}��]:�x�r�K��y}��0E���3L�a�B��4�wMKtcU7A����@�N�!���C��[�8�
�I�t��U����(���YjεY��5h����4@��Fta�Kƌ�.JA�#�����`tsǽPB�KZ�&�3~�*N��EE������T'<���r�C�gbU����>�+$�?߫��'괏��{���D'e�_kr7�ayM6�v�9k�#[��U������̟��q�ӛ��M<�6��2'����2�����g�0���0Ǣ������vW>�	X��n �@��ˣƞ���^��/�/����������,[�28���7 4O���/��(���V�+��:9s<�i�U$��.CY��xfJ����n^�$�I�q���{,SLM�D �v���%W*r0{�f{��`�x:���m��7�gx�����E���eXз��͹�����#��khS&��Yc��Ueh�'|-xmD;
�/^x=��H���5ۚY?µS� ���W �CFg���lҍ!dCH��}���M��=�]X��\Rk��x��r�:�pmvW/�e������[�u �����T�0�[-�V�f�ک.[qV��U���H�yv�P���7�bN۬�+�y�?�ٞ����1#kT�Wx�Ȳ�zVc\�l'�fSt�x"��0-���<���lmz�I�Q=@Վ%S���	v�w��;g��%N�ԯ�Y����Gڠ��V �qh�CF���07���4ҝb�����[��o"��)���ٽ ��=�V�fV�j,|Z�X>�������ץ,������k DU���u�(32ȯ�pC�&��50>ݡ�/
�����=X���H�7�ǯ/&V�}�����/ר�c';��];�c@o�0閬&�F�@/ �hʶzZ��I�Q�Hm��>�~���kZ�f��Z����+���|-]#`I:��+��R�,N���e��ɷ�c=N3����2�,��K�����= ��!����5��I4�2C�%��{����bT�"��5�4���D(��
��}����ҿ��t�x=���J�_q;vؚǩ�Ӑ����}c���W�	�ζe��m=�ҩb��Όj��}5ߋ��n�Wc�j��4t�U!)�qC��(�pDн���������p��;)���n����.��>��`t*y��J�A����]�C#��-��fU��a�ʗ���������Q��3dF��������} ��p�T�H3Z�t;�c�+��v�/	��y�������j��o�^P|�����,$��ʲ�OF����S�W�X9�N/�A�1C�=�b�:T�$��Ei��g�|�җ+uLo��Y������H��jyadF@�b��۰ K��f
.���\}n�c/ѻkxbt׾_�uM|��b0�N�i��"[rxI�o
rz?oAƟ�a=�o[~����q��B��æ��(/A����|[����E��ok�jWtrc-��i_�R��B�h�k�*�4K�!	��XLlnfx��-���~$���NV��?�'?�eEd�R2Hh�҄\k�Sw�p�ՋE���)y�F�����`T>sQ�ThV���L<���4Klg��#��[E+h־��� S)�+MeB�a>�\:�o�G]�Zk�CV���r���X��#���YX(w_��9S��������ː��gS $֜ƭ�}�c��`�7�����.N�ײP��,r(>ͻ"��?����� �4\̞nMֱ~Y
��y�)���>��ZjI_b~5F	���Cv6G�q�gh��t"�\|�%n>�8g|�yf�U!�P���_H���A��h�!���a晾���6:��$���]u�:Ea�@ˋD����u�m�����;�P-�6��܊:+Z�l�F��Z?3[#Oi8���0sE3Vb�S��ðq�&�1z�i�'1=dma�X��^[�=��r����~Y~h=R&6��<���u{���t�&O�粕��{1�00��e8'E��}'���ck��3���P'�5�3GC�l��j�'+u.ǅf���q��)͖1Q��3�Ga�`A%�Y�|�R��b�<h�H�7��+}5C���@W�QP�U���AG�Q"���(S8+Ni�� �^�M�y���}e0:����2Էο�������b������S�U���܅1��� 
������(�yG쨀�.Sd<y���D��e�N-��ځ�E"�PQKש]��bi>�8�PG�YB�+�kb���o�H��tC� | ��.���e��\�lY����=a{aӬ�� 'S�"X_��������[��Ѧ���ǀ2���r[�Bs���P2����sV��O�����J=cቑ�E��������L�?Hx����"��7`Φ~`;���&\(�� k�$�� R�ȿa+���[�]~�
.�U.I�bVzO���b;	 ���woL̜�NT3c��I��O�%�5z�d�J�obr�,�jJ���L���rҶS^����|�6�sX�{���w5f�<8Y6ׅ)��:I���ǯ(�f���F/�⃰�`����P�1��3��-��	қ- Q�|�2�U���Z����Oh�\�)�S���|������c����<!d���"��u$Ƴ�TS\�ˋ`3~�e{ o��M�*�@(�c�*��EwDN�f�?�)�#�ƅ��Q�zi�O�a�Y^*�Ӹct��h�� ��Gv"9Ӽ���;:0���*����.��O^�F�a����=^p�g�&�[������9��Q鲎��z~�Of}'ܓ�&_������?�n����H�$(�%� ű�Y���nɧ�z��f|G3�M8c��L���{8�p�7��`�Dq��u�k��T�󸀳���q���9$�4#f3	P�l�`�@�}W~� �y�Ҟ����4]�I����UX%#թԵҧ�i��y%J�a���/HCw�H\�)A4��b�����dٸ�=���/��LD-��+����ݝ��a�ƚ�t�4�"�(V�#to�$Lʌ�<� �/{ �F8��������ۨ�6+�GP1�A]K��O��ҏX�eXa�t�\̛s�j_\[dc+|�?	[W��Y��V�S���s��3K�A�y �����JZʔ���Ł�ߔ�;�L�|�S:t?�Rv�Bl �j��gY�%+a3��������.�2�_@k&oѧ���fh5�)�6����1c�p��AG^�h=� �<�<�+,+�>%ӵ���~��gl�jk4Tr�M�:�u��Di�M}ȴ�Vu�����@r�8K�+��w()h�<S�7P��a���	�?�?�R̰
��C����,�>2D�i�J�P�}Q�d$쾗[�EOЇ�5Z�L�%#�PB��[��b<�|	�Zf�0�a�S���!�,������F�.1C"�̡�f����LJ�����8��������F$��fd��������cC'T4�����������(g�Ixݚص[?�I��͵�ðdoF��	���`�M�H&xQ�x�w�s�����[��z��N��vj��{�N
��p�լiӵ�C1���m\��|����}�%�W5=�E���y��f!T�hN%cV�Em^_aJ]C1��
��%�����􀨏&Q72��jaP[��/z�hk�S���3�V���&�벊�*�J��O��d]߷ޚ��T�'7��� �g�z��͓4͎�͍�fT���9�4媐ݖY|�*�	�]�"/\�4�7j���N8~����>.W�x�`�#�W.�n��$�R�y�eg�>Ɇ3�=�:���э}�<}c�?�#��紑�Vቪ7=Z�$�h4EK!��aSf]�1?/�υ�l��$��QCW`��r�_�r����jP��L�Y���9��f�e�����#l�/������S�P���Iܱ�n	O4�,�U�ǚ����]#l��{������9{/.@f�Oj�e	�z���	�:j�p�7tݎ��]G��~���ar�>eS*k�,�]%�\��q9?��
	J�9,��l����@H9y)f1�e�c�Ͳf��ؐx:�e�֠�e�3�X�|��D`�P��^�{��Ql���f���~�����G�٭��;ԝ�kы�W�/�`9����#�C��Q���#�W�7P�m��)J�#z���N�۳$}{O �X��kU(��kV��v�b:E��\���}[�xD80+h�աq�kFh�> � �p{�$�	~|��h~���K�[�'	��<��v���3_�U�~'~�װ��)�R�y�40�%����d|w��8dP����ɛ9���U���Ӆ{����MG��8L�gp;�kx��G�9H+�����(ڑ))}�*�d�]�~ -��N��	�^|]� yE�{�,��	��@��\m��m�Bo���-@"��X���K���L4uiA�Kԑ�*�Ã�����HH)B��%��!!�k�F�%����qݸU��B��y���;:�:��|DHjs��W�T�立�"q������Ҝh^zd��Ýǯ�&��G,VZ�(�Hj̡Y��ó��f�NAw��d�@N6�<o�u���ݺF��;CH��;=�Tމ���n1�����0K�}�����!5>D�s�'��\.����mY;�;K����ڔ9{N�I�y��+�D"�i,i'YN�	D��R{�R ��y;#d��ڄ*PB{R����
IǎFJ�$�5;h/<����%/��>������9��M�ƬX��FCs�b��)�|��ܵ�����97Z6w����ā欼�"JX5�`,;*�y�
��'��#u�s�G�8��4�|�u�=�LR�"zF��;o��%�	�AB2%��d�'T�;�Ϝ�y��T�q�.�(y��ڀ�H6��@�~�5������7��5��[����rp��H���xS��t{(��\P�)��$�,�pf
�9�
�bP�=Vs]5���F,{�= &��$�sΔ� �0�iU��I_�G��C`�h��Ke��
����pkK{`�U)㣷����9Փ9C�z���B�-,³B�7xDj���$[�����e��6z��B��#����Y��V�������`�:�L���E��x�S;{��6y�(�<���#���f�SL��Q��_:Jm{�!#kC�U���Bf�<~ �Ϳ�~N9�ˇ�J���~GA|޺hi>���ƌ ��ͭ�[E����^gB�!�!_{!�����$;$ᨌ�ծhK�j�f���ժP��{�A	9fM��r��ɰ`��}�ᛙ���&<xb2��,�n�C��
�a��r&�On)�yQ�5��o ���HA��o\	�p���.�qit =�O�#�C~�T�
�ϯc����G���#�O8����yn D�@��8�ɓB��x` �d��
�ϯ ����)Y�HǞ�����p����U,�¥}P"�_�<�����W��L�)�w�Q �4�K���YC��x&+1��G�Ȕ�}�	���ʤ
��Ja�;��7|YHk�%Z��c�/���t���*�B���~=��#���Z�j�?����W�uc�br��M�Ǯ�Z��7�`���#�dxRu�L
C�Gy	�72�Bd�X��h�a��\F��%���X	�(9����T�n"֕�bf���5�`��)m!�zX~C��mK����A�BM��b��kk�m��bM��"t�R��E����jċђ���u�]謐a@���~�h>�5����}�����N/6;j�z�'	Ce�C�;щ�1����8���E���6i� ���k��|}����T'��'�r�j�<���&'�"����;�ea��c�V��E��!<��a�
?�Cz�P��Z����m�l
0�;�%/��_�Jnk(�F��;AjXn�cf��;�e��!Ĭ��7 �<�� ���7b`���O.�@�V2���*w$�.��S�ح?�L���}����\��N��U�/�!��D�7�e�FHAmn�N����@9˽ַ���("!Ԓ��/�eu"~������>���(���9�~�S��J���E��I��J�B#Ѓ����NV��P&�LE�:���瓾Y����Aſ���^����/�E��Z[����h,�OП�Q�H&MC�D �UD��U�'%�+V���ϊ}��|�m�+[�,�H��\��3��:^�r"!ұ_r�1����C�iB�y<����|�RgL���*����16W]c?�o����������ｂEk�)��?����[��=�6��d� O�f�=Y���}�7�}�q6���W* W��p�w�N Z�KtWU,���h�;��R4j��)��̬y�4�ܧ����D�c�����R~��:����+nGG��1b{D�Bi_�.�4�Z�����uh�V�':��=q��c/�x��J�ux��i��a���	@���l9�p��¬/!�N���oW�*D�|Xt��7;4�v��\���c�d����f@��j�֍�������q�\��o8�4�a9��MUw��-��=��=�U	7.-\���DJ�7����W�����"5Ƞ)ҝ����f�/���8[����~ן��"|��)\ɾ�����1�����r�_���=T֔>ȫt�#����{�h�f_N��M%��2�eC�[1�r�-�D���4e��ȢǊ������#%r�'J��;+��/Y�].t�"�#�'�
�Ov��$��̃��Md~�!)UbƼ�L�[��q>���/�Xj���,п��_26�-Q�WݣOzvq+�=�4��-!�ޕeS7}]����!�CQ�y$ߥj�@����˴�_�,hE�5|��f�(xd��p<��a�o�⺙L6kƙ�L'�I��Ag(g͉�R���@��b��M�@��f�]���Z&��^�Q-v�6��ݢ��A�;L��I[�8%Ca���	�yW���ќ�w9�	Us�y�CĞ$5����|q�t6��DG$@�ů�.H���J��>y� iQD�B��b��V�N/�ל���AQ�P�:��j\��1�ZU�<2���y��L��S������3z�rN���������8��}�'�Z�J{��e�TG�|�醁Z�����g ����]x����P!�����s
�)�4L�
*g�
�\)(Euh�|��H�cB���R�V�i�g	��ҋA��S{b� ����	h�}�ݭ���v��x�:pW^��n0�YvX�Ë�U#*�z�̕��N�Wv~@y�4����t�s_�[�MA���͵)�P�{]�
[|ۮ>��TbM��(�gRt�v�7�Y<���$gE��z��\�v��c'f]����CK�@쭔{y�����tq/�k����^n"l���R�g<�ڲ�x ��#ٹ��:��ô��q��6�P��X�Q�D�`���v��R��j˕PwU�ݖ�{�'����2s�Dܕp��r�?s�2"x�C�d��:a�*��x��<����A��F��.|r� ew	ا����C��Պ�����E��))Z�;X��y���U]�.0S�44��s;$ۙ�Z�����T�^0��Q,�S"�S&�������MӐCmn�1�'iu�aͰ-�.+:��s�k%<��b��V���8��ܨ�pb.�_O��|�ܧLj��:���x��H�CM+���f��eN�b�����u:g|��󃔕�ڼݐV��qS�Ď�j���^n~1���f��~��JCӊr2.l�3��3-%�I�6�E0HL�9Qw��MOh��;���	�YP}q�^���4�`��A*�-]�?�C��M����� �r餗�F"�؈�M�"ʸ&a0�oHS���K��q�j˒��j�_t��Ǘ�Q!��5Z�z�����MqΨq�8�L�3t�K��=ed����{����L\������A�Y������,�HΏvp斁��B�J�3N�鼙-�Ԥ�� d��lW���X���
��{Ks��q&�\��g���SS	]�N���ux.�M�fr�C����ZZrm����ъ,��ʔ!2�ո���F���4LL�>4@���m��z��Rƴ�I���ͨ���rT�K��������5��3��-H�v*�b��&�F���6�3��$BPEc5�V�݈�����;U�xG������-��Q�Y]}�+1���"����޷��𽵫�����z=+�R�7���i�	eU�|CO�"��Vݙ�bT�Q��('������a�Rø�t�̡��(��n���G��>S+��~������ۉ U�Qc{
��N�T@��@\����m%ء�����0XOUy	�����d?��\����9B
\�s��/�Ї<"�b~AuJ��D�WΏ"�W�ŕ2^o�|ڎ]��;��u��s�����`"�p7�ǳfh3w�V�_\�]��Q��z��o�k&���Ĺ�+!Y/����T�3	��F��h&��X�$|@�}���z��[���I�-"S�K�c�Po��U4�A3a~L�:�|\,Ē��-U�П��T�ʷ;8dA�y�a�7�x��,��d}��;��k�8�|m�܄���I��7�߯�D)H�U���Ho�^���A��'$�b�K���-��Xv�&Di�2Q��t{QUL1P��(Z�t�_�!�X���9�I���^���R��[�����C��3���C���f@�%༔c�+��b/mrh+v�oBBC��vf�u~�w�_V��MJ�:���.o��m]['c�i�6;�S"��aW��	��e*_;E�A}N��3��U[�oJ�ݘ�T�?��Y�"��5�wk.,�X���w��Y� '�Nlyw�����S�ӿ
M:%����M�<Dm�����n.S���I^�P���H���yt��n|�0�3w�J������kU��e�F:�0�S|2��X�7��J������Xvf�[?n�⹱����"�̏�0��@VĹ��OP��C�x��Az����A\���D4]l'[[��O�`�jJ��T�;:�[Z �?\t�UJ����E�#��B�z�B@�2�Ry�oл����~0f���T46H�`D�݁����Q�,$��a=����G<���0�O�kf�7����E���[�F��'G�����%���b �;����p��m@�!��d	��ǜ8@���j80]'8WH��V��jC#�o� �d�S�FQx�����-��aK�h�P���^���}"!S����Z��kѰ�L�x'O:�ן��d��m*ގ�}e[�}�P�w@Ե�@-'h+U������O��,�!�
�� ��{2�����@�&GM�WR9X�u��8Ѝ����V��q&	��f[m;�@��?@9�pS:�z}'і�9�T��fvp���a���|� ����GZ��>��_IR@x��j��8ˆ���ӵ���5�V��d9�&�Ť|׆�F�b̽�����H�}uh@�y!=O�����0a��k@B0:�YN�+���P��J�%#�1ڼ�ru4aG-��CAA<E�����^�褟A�����5&�5Ě��{@R��Rx���$;�3L{�$!��p��ܲV�{�:�fPRE�|�\�ٷq�A�c���W��X�Zƿz�N1��'_�J|�M4�161�
�Gf�z|�����o��J����4mu���zm�֢��������a�)p��Z��R����f�.�R7#Ѩ�0�}KS��zXd�����0B�0��2�B:��g����Y}�A+�6:M��WFB�qؑ�A�X�>��\�r3���#��K2��C���!�����������Q6k6�ZxV���kA�!�twE�W����z����=��5i�q���A5 ����t�-�8