��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK���mkݛq�K� xwC��f*CU+`�>�zkS}>�����{���K3�&�4�N�����Nؤ	$̂lUPo��t�-ME�U��j�Ì/����$��_s*���j�^��<��
�ZJ�S����C�N��,�J�e��$,%�Z���i�>�B�i�1~X*�P�}�.W95�f1�t�~�)��³O`��P�d�n�������P+�;���tFP���yr��f:ɽ�N��A��s%�Kc���Wq�5��6�`�{@.(GkC�7��aFgЄ�ׅ��+�b5/�{�c�Я��:c�<۳����]
�~��܌����G,s��۔�ag�H�Y,d���>^�H��:�ل�40ٝ	��#�<CQ�����h�2֒l���;�D���a�����ރ�簲{:��l'tJ��~2�w9>��3����m�F�?�8����}
�
���'P�\���J��(u=���~�$v5�ņ���5��:)�/���$�{�M-��Ʀ���n���_i�S}����a&��y��3�_��-��ӹdge��ȷ�D�\C���!�]�Rk������"qf�pN�N0�ǝοg�}��v��c_�fc-�`a.�CUw��l�R��?+,�WJ��tFY���dG���gH�:J��".�؞u����Q���u�OY�Iy\�����G����4Bgj�5�.��#},�_���#��8�g�j���?�zA��,ά�.~����g&Gj
�l�k���8�������q�Dg�rv횡7��/�2�Z��&0�PU�Dc$���õ�ER���"G��a�;���b]
����4j� H��[���1-N��񌳃����x��&�͇��0�f�e4[�x��G@$>N���R3^%N�=��^��BzV[��o���kL ]fW�����N�'f�l����
J�uc(:k���Ze���o��q
7�����W�+�����8R ��Um�c��*�Y�tš���q�&[�xd�����R��yc8���k�#�	~�9ۯ��`�{��72 y����}<��K/:��5-Ź5.��T�@U�ʫM��M���V��
��֎7�Z/H^�M{��ݥ;�k�4��Ԓ�w
���+SIϦ|X�g�~V�;����s�)��MkJ�&X.��n˥�|  ��z9�_����	�,���jK����݉�<k%�41�_o�Fy�3���?��Ƣ�X�m+�h�f�����R�� ��ڰKeZ���$��Ǻ��I����˭}N�bs�V�qߺS��+�>*�
 =���\�l�o��T$��v*{5$5�b���I���l�ra]��v�c~GSS':Ox�)h��>��dZ�,S�rj�8
0�	8�b�ɳ�V��i�Tv(�K���rB�`q��mo�|�g5�A��g�6��܅>�M��B��J�P�jW�˪�R�[�I$Jc����Q<�J�S��]B(�����U�Q+I�N����w
�%>o��T��|����`�!8ɖ��3'��S����[u��X�	_�u��d;�7���� ����e᲻��Z�ems,����=R�i��[�d��D��"8��@ʆ-ݲ*\���30�d�c�A�	l�D ����R���ӯ��3TL�L�]��:+�Xu %��|� 3�SuY^�Ňq���7��CCΌ&pRa�Op�g��ES��н�2QWK�~��\>:Ln7�̈� 9tW���e�ۨ;^%���O%�85�QӞZU�S�deT�s�6�����7қPV��%��%)Xs�t��:m*yQL�*����WLB)|���˶����7m��y �)s_C�i��Gȫ�i�]uCdH1MX�xP�9�N4	=�b��u����=|�x��q��U_I�j��UvY4zj�)��{�@��!�#i\�3�`s+B�
G�V��g~ �:���zX����ET���1�:�N�BJ��D�?� ���˖�ha����J��l?���9zUn��ѣ�J�dsX�-�4؋_�G���z�"Hx�O�� K�R�Ң V	 ��x*�g�+�:A�6roǪ�S���(=��~[�����
8I���;�Ӑ��w(�$�a�#�z�|�U��S�P}���Sjy��'A�H-�Uχ8�E��q�|y���;�	��F%y����Y"�-t6�gw�5FK� ���ǋo�n#�7�_#|_(IK�Q�
v� �-��]����͙ *f�������Ã�Ժ�Y�U"�}O|]���I��\h��܊+$�Ŧ�+��v���H�窯������~���N� )���!V?����&��,\n��}���Uo����v+����k�&@<�qgx_<G�9��A�.�y�����y���y�}O��B�$�.��n-t �)����^�$)!
pR��d���Ѽ����'R�lP�"[����,��lKL�.�x����.�M�V���dX-�E8]�#��{�:d����4;z� �����O�+\��G��Όyڼ_��2~a]��vz�R����<��y�y�k�J{��Ǎ���d\����<`9�|����Z ��i�ge3��e�����~5)�B���-��sԎ.D�g��%<������p���f�Y��7+;y�@�-�:���iוE�%��w�ץ�.u4��1��xm6�P?ePߘ��ꤺ�fG)!�V3΢}�0J��y����j����@���K1ߧ53�M @V;�'��BhOW�d����K�~�*��	���%ZO�ؾ�u���n/g,�PP��ʞF� k�3P��t?����-ͻ�������΁*�|w�˅�sHԷZV%����HpzAEᘸcu�S���o��>h���Ky��o�i�QQ�\�X���`p�=�	����LK*��ѻ[�=�RCX�X{�8�Өx��6����|���1a�	�	S�f��P��f��-޴�F�&��n.�7֒Pܞ���5��$���[U"˧|NG �T�����u��Va��l� &��D�zXV ڀq�+����ds�B) �=6���f���� J�Ql_bR��4�U��K|�M
� 墕��.<�֢�Ǥ��X��X�ZsR�مF8��7���D:���̡��T�������e��3��Q�ЋED,|�B��,=���u� �3R&|��X�x}mR^�83ywK�RStϩ���A@������u���i�Ga���y(�7�<����	��!�E�#�ׂ���/�X�?A��Y0 �w�΃�HG?��(ӌɖOY_�ڇv��D�!w&�)�8�)K/�B�N[���0�������8��VAA��Λ��&ONl��"|Sd�f������,HSaLSdC5��	ie�Bz���xp����`Q�K\����
�����H$F�<��\<�s0bv}cC��(z��p���1��%�ro�U1Mc�Z�?�u�mp�D��6�vhա��$���YE�Ҏ�<_V�V�e`:ș4V��UM����ց��ݭ�O�+��;?a���F�U�x*� ܜR��Z҆W'��|���tm��$�Jo"��NF�A!t�Ƹ���k-���cŇ����z���������:�ĥ�j���h;�}�NRZ� ��,�S2��z��&Vɽ��?�O�z?��Z\X�LzgA��-��˓2�U�,�z��?k�6��YF����mh�E���x�6;���#*a�qlz��I��;�G-`�چ��r���r`L�����׊O�TV�Y�;0�����aPo�{A(&�h�)��3�	��o�j�X#�O���"հWŌ�.��	���<��g�-�̏�Z�Q�z6�M'nZ�9z�$����*�N��L��)���~�v�J	�P���Ը�>O�=7�&Z"�ow\[�n*{��p�l��u�D"1ZcOܝ�64-;��� o'�6�z]nMk�u|M�%���m0������D�IGv.勱��;���6��~V�#_��*�-s&�i")hk:�o�r.ngi��̦'Yp+Zvɫ����O|�^�<Ś�Nis�=`�,J ��R�!hX.�#w�cлǥ;A��&�я��V�_�'Z��Z�X�n7쪩��������_b�o�7���]t{�8�:���!g �9��rB8y��ч�Ted�Z���B~�,������">����9�T%6��=�|g�d|��ъ4V�/���^Nx���3��N1�"֎vU�[+,#�fO�Ky�梱�i? �%��b�i0�b�6�����T��p�J:�U6мU�D�Ն��+PT��`�U����A��"�}�����AVt��᥎G65�Oک$a�)J�?xL�(������O8��V�s�ǒ����lDi��;I僒�P���x��84�����ԦQ�gٝ��%���81�0:�3��FrR\�+Zz�>�|��R��$��]�[�~��/7��.�j�U�&{�H������bQk!y�}��OH�vhd*;�FVC[�St�,/RDX �>�;���|kʫ�C�!*axV��|�V#w�X^E�R�DKW6xNMl�#VHu�Q� ж�ݭD^jÇ�=�ʀ�����aqj54�(,<K��)�����X$Q��=�K��H" -�.\tL�8����[?�	�1�|İz�%���G3��oD��K�H�/�[�M����؈Si�8:�SO������� ����M���s���ׄ�Xk����4iO$K����q��^��8`���"1�b!�qn�=�y�ǻZ,�"�?P�ГmI�7{���e,ϐ�+���?�d{X���u���ϵ!#������G�èS���5#|�/���Ϥ�ZD3��!�.c�����Q��?�.�a?2��^��fӫ��Chd�aP_�2l|�86yL+U�����4):�{��<r.���T��M�p��gl/x�,WΙ� E�Z&�Ft�I0�M�e*�_��ܤ?�Ў�k<���B��Tcؖ(Y���a�%ʺ�D�h��T�'��n�.TB֝3QX*T��3%�6���Z;�e�6�M[#X`��h�&��g��ߋl�sI���5�V���p/�=`J��&%����'�$��T	
pc�4�@�r����C<Y�_������aٍ�7ù10=��B��HrU��k}�72�DܳD�b�*ת��Y���3�:�wq�Y"��p�M�#3GsF'�3��Z��"W�{In�r�����k%�o~$Cuy���7(G`zO�|�w~���H�/���A#�=�U�|ἦ���_Pw�G�_�WN�zط��b	Ku@bF��<��@�? fj�o�����Y &�������~��O>����̗gi` �%��C��*�n-�cN��b�5��G�̊�Sf�c(Jm<Ml�q#$wU;�#zl��K6��󒞀h�$�W�"/�ob��jE2��?q<X:.��og�e��JH��J�a��4!,�F^X��]�m��$����a���2��q��/uGZ�R�S���Ԛ�s&�� ��a��K�"ӎ�4i9��� �\�'נT��=}��#�[��1hFu���g���sS�m�ޥ�LP1S3i:֐r�w��o�*��=�����?��1A��/���!3�м�1����\�nܒeR��wӴ��Ԇ7��,�Kd,���@��d�Y!!\z�Y��c�po�׎+?y���%���Ż�v���t����-L[d:�@Ldy��j��=z7�k�H?��> �[ET���e�!m��m_�I.k���nI���'��ï�;r4���7u�V+~���"# �I�V	��N��ۺ�x��ŖT�~0�6�o�?߳zY��.��~Ǌ��fߌ�v�Zn��Ɉ��y��_  _�a�RuH ���ݟ�M�k,�I=�'g��3���8.J��u�n��ʝ;D����y&����.@hg�w�:,��A��y�&�x�&\�i��:s��qOn2m��QE/Y����o�0O�b[��H�P���0q� 
�Z;�ZT�Ý�"I��=/���z�#�}X$/[�./V�X�*G��g��A%�m*�r�+2�2L�uRO\({e������X��i�Q �\ ��b���D���.7���AF�Q�4��1� �޵d��|�|�t&*�Ҷ�� �,�e��<(�H�G�@"�l� �6�Qr�k� :7�D
�1W�/�
^��\�����*�e��z�T;�K�u��#?���P�@)Cm�������@1Z�B3�d>q�������3�"
;���Ъ�h���/����>�����|[̠�N���^j���Ύ���SO1��wPOg	�0Õ❗��F��VD�.ZM�3M�T(����D��E�KR4�%^�
-V@����g��3��H5[�_r�Fm-\*���tݷ	��s�`���9����)%��(us�:ȸ�Wpp�\u/r�-A��m+<�tƿxSIZ���p��'�-����T���e�����a���7��������̐�^���@��&��������0��A\��!���F[VWvY�P�쇘���؆��k��-w�6d�&'f#�/��UX��Z�ii0�������N��D�I���y
���,.
��d����Tp�y�b�T��c�wV��d�����-Q� V�f�ԿC�ɉ��f�-���r��|���u7[���w���2ȿ��
� ��H/�ɋ�M�}<��pEHF�|�r�H<i(<lϨ�'A�����k��~���<�AG�H��7�e�7\ل�t*=�5vts�}X�^�'\�2�3fv6}�?���=d�Gr4�EgGڦ�IJ� ��'�	�p�臶E��87l ������*��7����N�l��[�k]�2gK�+,�%��x��v_|�1'���?S��_�� D:?��v�T.�pa0oL^���Rv��F�b=B�q�^�+�#�յ��nK���]& �v܎^��:q�ʋ5S��W��oy`n4��-\RX)NR �O���p@@}�h��� �>n,�V�q�A|H�������Dl�!*?�w��ߓt(�]�>��|�4����T(�@����y�����:���w��V|����O�OXEr7~�;����~3��z�I��0O��*:���"�	~��{�]�� �=�\��u�zk��DF�pK|��tǱ1�n�N��/v$JKʭ�n��o��(,�
�]*��k�c��o�J�S4k�
S����>w�t�$�~�MԻ�L�BR��d��-�|��1�$_n)	30�}�k��!�+�f�0�}f��u�WC��
���,e��K{b�i�2�SPt���.�r�)B��>���G���
�iԔ|):�b�$*v��A���Ѳ��>��(�E��9z�`���?Q,3k;����*�w