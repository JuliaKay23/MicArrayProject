// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:16 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WDU+4yI8Vr4yqxJSszoTPunRThUA7xiBbp92AbwwJdV3gcLbFpmM/+/cJ1hw16zP
geF4ixkBulA9BvW7hKPQUpDeasNOxITNLc/5g2FFGTw4yY0R++HQnYUpr8bdUyy5
18NUrIxOUFv//HsEqFlVKskGt647pIORuUHTng8J36U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2064)
T8KELgqAFlsubdCM40Cb1rliMNY0OruOQ2TJ3wcZfwicQSCk2+1SK/R9ZCMzwCSo
imvIpmAD3+5obLi6K9SJUrcLXuockIobQ+4fqETGUe/6fHbimTl2vQqiyZNkwB2t
KIwXnrT7gX6uOmk9ljU/CC0LxxsqHDM9flIP8fE2yNQigZrNOe2tdr9PFzLYkZuJ
xvP43BxLg0wdHVdZ5Fa5xVKjIsk5/x4lW6B0kHWeaf0zjDyiVUI2wTZTEnvyVe7m
PcPiTfU2xeY9qbQcO0AMa1FMl9i9BX7AOClB7aQqmkECaWJctUJFE8n1FrWa7NkE
6u5KJeu7Sv8USUl193VzkOFO/JucQ9/YZdJ2pDRODspqmt2ng11sBQyXCzjUgBoe
DcWu7fjpvOAzTNPyFGqCIWSBtBqfRFQNbgWJ1O5D2juLp5DLoNtTPqq5bRQtM3VH
v6+PZaWPYynlZpb4kHJ/X9lQsfzmGwyvhdiP2H2fY/lVuF9LdgAAjNn+HfnCoahN
EujZEqS155Tpeydr6fAn7iU+i3opaGw0JseAH6xiqmfju5WKjgJ2VLcjbFbP5XFz
K6X+yRaz0/cg1G60iKUz5S7LasIVWZ2O0r9Prgv2wwjbh+/0/ebe5CMaiNjnZZn8
1Cq0ySQ3qozSfv3M7F0L6lLOwxpsHPm8htfjvIMj7qYw9nJh/EKY+/Kykjob3+Fl
hMmT0GUE1S94PIjrYXP4Wji87HfpxxUgpnMf3GkGhmxg3kIL4ubaI/ecbC7h+PWs
za9eb9Q4OWFdtbhftcuPpJaJG9TUZjp3rV8rwpLFQwOmYkpjBQbJpTHUP/FTSbyz
ngUiusu7f2sTh1pUUD7dZJ+L7K8Z5HHb8X37dTnxvlVhGgMcJyqRoSRdALMX7ly0
vaXVp4rIUl+2Ql0KFABU9fqUKWGdGW5c3QYFrGNOWloDrZ07+gtF1s1VDaaMhJSz
MVHUQkzmRsNEW+zq+4AXrftUZ1DBJ3utRqtDj4ETlZxVys7xluhw5aUS9lhpVIeX
c2tv+dRovTwKd9prBfhhdBCMjJWKWE6Iju9gzKm1N6msr66FXHbqUV3+YCVzdIAH
rk6x3IPgE7Hj8TXA/UcoiYTH1iGHH8cq8lkMFafF9AXvQM6z7yGxrLqxTntprWtq
oU0r2KQAY5cbJcUFQtodL7c3wLcHxZxfKsFdW0Rez3MijgYYlavtDk0SXsPvVbM2
f7EXxkeWtwi54+h5NvV5SMFANvMx1AxzQkGKi0PcW+Z2omMo8JwhnUZjh6u+xg6B
9y5uZiFJ8V8YBcdr3csWA60qCTEMsHLC468x9vsXUuubvYw+g3y8rPi8Qu6e81Yr
5jEnJ30mVrFbpIPMHkcyiQmSzWYuwYMHEu0eq1S3xGLv786Hf73/n4hItisGjba5
BcKXRUduaddU4j4X9vO67+xyG1jA+ar8zGGtdiyFp/RDKYlxJZ4Q14pKWBZbjRqo
PqV4Wq/YX0hcHD5M+CmUwF+4CaZUG57b/e8vTvmqwtoedRGdN46ght1gZYGdqLFC
qF46cfxpuUGyrK6wpd4eQrFQNkTgJ9bgq8CCZAeQbxcsndBP5GyK8+G9LQADnyl3
wz3S7Vz8f3xh/XlTbQdLGkXnbF/lrde+9r9k6aIdmJ8W1mWIIzUu84UbrvqGA6OH
iXmQyyHDXQeTzWc1hfQqjCXQT0qyEdsudCfgJ1518aoRttkmak2m7hrz/TPFh4uB
QL0KS1Z4EnOTRzdGnUcZsW27zEtKbF4tXFVcJ3Jo4q6bJ72qdWaTC84M29Fe1R6q
LKy4+OuB8d+r9/LgXkYhiUpN67ZbPngOlpB7km6i2U7T5ccoKGtgGw/QJKceD41S
StdxZtB3Yj/kGSoItV/PP2Ip8MTYWfCA02cVuaVOtkGJzB2GO9OV3qLZyNx0CV0y
F6uplj4kusI25s+91Z19xW0EKukKXsTcSndk1jco1AQ08yXREmHXuDPcXQeNyKjT
0MIpSkWrjhWacgvPMggvcEfAz1zWAERr9kPBZDerBpPdUtaGQFuwojSmqelGx152
oJsQfSawTaC19mCSiYL1x39V43i947ckkZ477zEQbh+T899dddv2yGw4Vt3prdwv
pe8jIOtXy/UvvkUbg431o6kewqQq/g2+yzxFCqSnCq/JtPbO/I/19UsbeJUvkGkA
JWReuiSd7dXbkZ+A7Vy6FLJlI+v8UJWmHuhZv0qBfRbXUWBgAHg+sHkEYLp/eRrN
I99JboyPyd56sxZOVyfaXfHUtvdqqtvMJsY7rBcBzmhYqWWU84PMoRwP/F+ZELkD
LpMonA2TSKqsfDRW9itAGHGu0P2/nvYkfpcgFqEdOycbfEHZn9obs+3TEC82Kqo0
PF9nD3syODO7fP228a4+R2YGlLtupfiq8RKyrLiDU/G5z+VVqydryzB9oILrlPIq
57WklcRPV4EjCTSBqzMDiE7FdWzssom/JoOFzmnJ/4tikjX2qKDN3abSVshNjvwH
xxaoxcBejXcrZN649kyMXRfppTNlZ2A3r6RuNsA1rMx/QqxCZhqKHYSXXVWy6jKu
3E7pn7hJ3s3lo620ty6YZkFZSKKJnRmeMuAZxB+mMHI2SOS0WDvkrD26OZulUwfB
zDc8b4nmmRsTajch2lgEpl6RFcxrmq9qr5ab2Mngo15gPAiAR2n83iReS5n6L9q0
FoW5giakYO04hkEWJNx76wQXx/4gBbU3sUzMC5IEJXA6wIu6GHdDSvNdYYe74tid
`pragma protect end_protected
