// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:16 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hLZrHdzu0rhGmIiLrp8gesJNhIdEd6lDB/vqV/QpgRxnNjPcj1umGxOU1iD6ND1k
NPCxAHMVpw0Tw2MjXCLURF50W3/k79GRu4YOFQUuB66gKdLD4iU92jfC6xKfRT1S
thH7EocnkqPkyLnRWv6m9BBmeIl0I1gvZmpxF4v8f5g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
KCFO0ppJ+EKPTxR4pjudIpGHlCDBhl6itmBRpVgggFMMwcAkiZvCadKMoxA/CqB8
PfdnFrB338QUSe4HllrLcwaBJ5m1uBu9BTjeu5VW9rQxoYAK0RT+C/1A/S88yaIG
splI4tL8XBTBUTmewWf05atfg5AFzn9TYfgKX2OwwDoWddLJhxe53vBZ4C0I6wW3
71NJD1PN+D2OTBnyB4+EhNCCzCkwpjs6RunE18QjD8zEhz+LqhpJ1zzOR7J+XtQo
f3QRcEqeN7CtrKZ9/DW7WcfiqEr3l7IXJNw00kM8+z996RrqSRAiSOa84QpyyckP
ZSTd9BYbG2yXsuO+tR4p2YAUWecXAGfjcbVFgVeXMob7DFoqfMEzdKy8Vd8XygDZ
e6sZ9N9kuWe0WvwErB2UosuKxdMiAuq5uVMWV9pZsV0QJVoFcyuO178iUcoN2pJW
6xX5IwshbhsacAufV4fY3mUJ8xR933Fl6814GBkvNoRUQS4tuEWI3Hqnz7Z5Pu7b
LgRrI9mwkPvyQnQmqm4vwjnW3Cvo+L3cbHZjQN//Bi9yDoJkfaBkmY1WW9hvsglX
fcTCV5h9aMAm6N93uz8YFUKc4fHWfdNQgTDrsRlqqrb022oXZ3sh2s5wteoUuzve
9K10IugHtWmanFSUv/1tKhgVkJlqk22CRFmBezZGoCD6GvuBLVIdw3lPjBLWNY6j
MAfx3zD7IvcgaEiVYhhnjILxTgpDK6bfrp7Q3e9YlRops2FXgk0jExTKfGPm6VM8
Z3XA2BDDYpBpgDG3UCiwyoX+gEGDJ/DUKKIioMPBOZNrj+6jqHc5Mk6AREJ2tbvB
FbNeSdsnE8KTEflg/FgoWRCNE141ekPiNuGV+AYv8CMRCngPb+f4BcxrlABX46xg
Es907xIRlg3ISwfAqqwJJ/Hs0ovhc3a/e8jnfMkZZXbEB/14aI/WOLXZmDE2w7JV
Gj3OtYkyfVBLRCShETVrp8cL3Iuzl4iEg6mN70ri4c5T7hG1J/d4MU4BiLxzdFrg
Kfzq6SI6tnk48VihFSVwFyv1x6bmWcrpEbiKhQ9eNa27U0Uej0IrmxH2s+yqZstu
4l9/fqjcFp7gKq9YP55KpxjywJSMCxqG+fshqJKXuRWF+RlTVywW6PkQLqvusrrh
7SXDnwO3x0O2LMc7PCXZ7Ly1POtdq8yPdmoPz85/FKIVqqO5RQmGpQ55TxpEKncg
U5y9fOo61kgIaSeB3K/68vmDp5yIFMnlLQ3WC2yCQ3Bx3HGKmGdohF/hf2HWUeF7
8Z9dwIliSHCYXnXRUxmVriOz3mtzBNMk55TnKG6SUgt2CO23hMM+9wZE76QVnDLg
b23TrbNzdsldO5kXRe1k51hZtOJxD0r5oGVSw6QVxE78osT6M7G2Vq/ntE/3FSIw
058qyRmaWCVaGMv/khYAyrtZ9AIivXTQC6EpEZM25SUkdSMyVZyqGSLZEhSRhgf0
Yx7mg4tcUI4fbGLYwjNijwtVJwaUxsID+3Z//WFI403dhsZZMgCDEOB1iyIqdANm
3q8Q/PUdaQH4MjqHPC0Jlr9TgQrH/WI8ZFKCz4ML9bDJ3cV9zaBnNhPpghZDWlQi
xkIy6joAV4BNSlN8TWSnw3eQikF+GL+isjtt9xLaTyepjSgKUgkXlsXF1Iyt5aX3
EKHDhdlEiYrAcdUn5w+AyO1C6GQNsKZi5/sr/xjPnYnA12fC6AXHCdIIl9azZoUK
EElye0bDbtKWZBajTHR4ZDAEQNfwJtAfNJkfwwzMOuAkwzCq/aqNWXrbAoIP9txP
W2SQV1uPwNJwik8b1fE98rAFtpgPR4o8zu8UE+etg/NLUJ38UkqDMxTkRh4F4qDJ
ib9Q2VITqq9/3re2c4slttTIjufwmCOkHsYoqv936eEQR7nBvf1e2avT2006b4/X
92MbFjlh65X1jRxqJiTK5R+QHYvMoqMQ2w6wwhTjnpeaYUH/IAWOy7EQ+lI2XzYT
Mw+xQK0WrpSBRUmHN6AgXC3oY+9zA5qCz9hAQCsjFK3F7pSSNxGGJMAEj0j3iZN9
/dop4SNOCxmlI+LuCnOZho11Pa3o1XV7C8J6EvVUei4QM8dMjc2mmVSJe1A3E2Og
1m9x3GKYQxx5tgoxJBKMxUYkVO+XlOQpiBlCkdXeW3LipEoB4oW+A+wg6rUr1s76
cdedjiugt5e1AqmFr1bNv7WtxwxoUXcp3s8Mk+AE3fu0LPRdSKpjNRz/sRUle8bX
eI9AOZvdVpB1sqjr4NPNg9lmgnxAedJA5KQWgp+GoVrL+goJDhpdqit0/AznJ7ij
c+jmNn+AEHX2Eipvhay9Pj4Xo6qw2pqnPq1MWkQ13qA39yIeWqQejY+0hCzOATAg
8u66Dq9lv2U0McaxRmZgjG3986YdWBXDFEualvxpAR4wAJKJFxP+OjqhuTLT4/tp
lGN91PiMB+zlFf0LMQsz/b9Y0OdxGl8sTd7NlOWtWz0/hXIZDWa/8/3EbhOnjCdY
AS8g5tCH034HBD7bvxznsrZyMW3kBynlRIfXfPbphvc5YMhhW64NJTifYkq5C8aS
4SWUZ3YmqtbS0oY3wBwSAL1BKrZDuWdiUiQ8pmjFs/mAszDG+gDH4b4ayOb+Hcq8
s1z37+keihVCH5uRKkDWiU6YYCe5vBI9zw3XzMC8sJblZd+zjIOXGIuZdXhqU8Ll
3IFsDSVQBJBGQZlZMrVlUSaLoXjGFcW0B01RKDzPZsmwPEdfBL53JbNFHTNsx6+s
Bld/CwdharxkrIHeOhHP24DC0xs29MswdYZ0clTonZT+1SgQbHNATUkNlKlAk4V2
UYxyTMmSE+JPMAAh9FPiKH6CSR4GhhqTeOsx9koL0JmWsmROhWbz4I6TQNppsDti
atoPI1F+JTreO9QBrWk5h6+Gbgf31TCopnjKBb/V+jCqdgPB5hWCmLT7Wkvhgvlq
TGz4vjPJe4hJdGveJ/1GQ5jiWo5aM8UvLJPrHyd9MgLisLJH1aY00OJHUrb3xLzm
bzy0MUtUnbV8Dkje0FWUM4Ikf9E0tw5RRlT1iwJUOSj8EsrK9dD8458kzHWl0Dy7
u8K4YQHz3+TV+rnJgoAD15TqxnAqCe4IzB8emdZVRGx74zTrGMSDhD/eUPk+prx7
LUgMNiPww17UxP6a39soD3fYSEaUYdM7Ltu7aUMFtLAZNCk9PcWdkfRVtXaX0YnT
CcFDPcqI5Z3fT0A6i3ej1YMkhqGg+W0yrRMKkwLCzwXdsg2OBPljMyxAtk7aGyU3
CzCGNkiuLDk+KD9ACsZh5Zf/EfrOOfeZJiJHNPplQPdCLuEl0JNz/wqIH4xwJiDr
4I+QwqmWjdmcLnR0eN9eioi4R8HC+gchKNqJuTrkBtyMz69NIu9P1iSGhFuVmaYz
57fTwXXYoiuzlE5vh35tCZUaEljtuUyZ40YqpWtQqW0PKmDQ2qkYyzooQE8dU9ox
ZqlJqy5rRZOzshsrENhXwC94EPSvG7/RHDBfsgOYPkTuqVUonXJiMgA9qoqK5aWq
mi2hZIrlDjJueC85FisGOs4BiwlLhCTZDTY8Mvstob5QBUpaaHeDNcYS3/GGcbO/
QVsAf3r/OZasxVUt/orsBfliLixOlrwaaQwAMfpcw8ihHLPr+oSVn510LcMiKne3
UoNsjOSD8FlaiG41XSlRBckjYfHTltx6itIRxFtjgnlHFhwUioBNSLvudQ/rUMpR
iJa6p+URG1QD6re4B09UELhevFZHwVL8dG+T82x0IWLCFhZmbEKAl3rYiNCfMlx2
X4u7G9g83BhjDCgurDjX6jWKdz9Bg3/fSdq535xKz1E4nZIOeWF7AKWbURSpaUyr
5a+tSkHF+tmWL+4TdF8XT7XPqQ1TL3e1r47Frn4wc7itpEb6UWAqxqALL2sX2LD1
DSmmj3gTe/DOMiwNCaAvKFds5o9nDV53AiEXiDyb5k11QHGlJ8PgROr1YeQrVTYE
QBsXaDBTGll9kMtqIjyx2nCGpPb0zt/EN6m5z4jdNSLD4mUnQ1DIk4uhhKZE/nMb
3DxTKeqp6s7fs8bzxMoCxQ==
`pragma protect end_protected
