��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V{a�p��H����.T}DM ������|�輛����*�
 e��k�vn�e�WY�v��y6�^KZ�� ]L��(~��p���\��M��R�Y��(�h(0��!�������h�b]�6�������O�M��+�	m�F����1�8Z�p
A
Z��q �ya�9_�q����ԕ�����X
���<Q���pb����#V�D'��P�[w��s�-s�"6�/+2X%�`���	���돐I\���Fc�3�@�!j�@ԨA�)��G�\�w݃6R��O�]�f�=�oQ�~P�]�e >�-�yRw��`�#n=TI�/s��,�|3' |�zQq�~�@T���z{w�W�]�� �Z/3�o�c������l\�|\C�eӥX� &T/���C0�ae�U����J����{2�������d�O��j�`���E=���
z�{����vEP���k)�-,���#;Rr�y,ԝ�L<��}��c�L�l)y�.��6����{��ﳌlG��J,�{Ɲ��S�1�%RAl��օ!�d�j1�FZ�E��^�t�G���h$�#��#�яq�M��d&{8�ᐐ*>��ߐ\ZXU������hUǋA�.��f�A��=�f�"�B��ݏ�Q۱fY��ü,�_G0"�jT���v�
("��~˷��fK�4�s��*^!��fA��7�q��wU�]�"��q%:媩� �t[`6'���0b?砨�UxMi�&'V/��8M�9�Q+�| F��D���p�k�o�XU�#��˽%%0m�4�~���Y�&��н��1��֖�$u@���ZX� �By����a���nT�_�Z'vbs�� ���M-fߢ0�1���_{ ,E����n��R��aǮ�KZa4��a� �[	�(�0�]Qnm<��F����ď�U��qg�n�D}¾j���L���ODV�i�H4ҳ����赠���.�����an����gc`��V�U�}� �����m)t�28���*�(X��;Q��1��:%�o Z�9ۨ�N�o��3|��F'?�e��^����W���8U}=adv���&{��aTEN0����=l�z'<�%ZBZ�J�E0��v���C�^P8��H� �Lo�1�=��������s�_��209P�I�{F�h���ܶB!��w�gF��&��t_�6�q��*�����Gu7��RT�hCoI/tIrw�Eu/��	�� �no���NT����"[y�P�vȫ����D��W�Dr�4h"��4M��5�4Ģ�@�头z��EGgNT~��3�9�ĝ��V>����XC�s�/F�j\�zP���Dj;d�>���C�5�=M�uN/��F����5�q��]�6��AW�W�K$������cˋd7��B�p~s7fJHo]�#���f��dȋ�F���g�h�,/J�A�:~JVQ��� �`)�z�������Z�Ţ�'�����e�W�ӂE�ZǴx;sQ�e��$�/z;5.E�f�0	��]��O7}����p>���<�����6:���)�����Vq�ܗQ�
�q���D�TF{k0��x�)@	�,lJg ��#���D�[H�7��u-�j�{��&�j�*S��:
:q��µu�����g���k�R�Q��~��a���n���A����z�1�H�n�=My�H���^%�h@ 2=&���$���[C�v��t&�^ 9�S��*�<.�W��s�j\qxFF����A���9��jL6�����#du�哲�2&�Ƣ�i���q�I����v�+Rl3�aRͧ�n/Ȗ�vz���h̶��a��{���	��(5���y�R�{��ۙ���s'�6��N��6(8��A.���a��Z���B�E7����uQƪ��{YP=���Po�)X]^rq۾גb~T ,��+κ$����s�Q��Lm|�U�\Ą�U3��i�;�)��Ⱦx� �Tu~���z7�ߎ