// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
GmvXRWJB4VmPgN6k4kmwS60O6+LWQD0aFphgpRQ7z1XjDamiOygY59Dn5Mo4WCPfs2xG/qjuMORB
I6Cw76n0BXSclyROooq868u6g1qgh5hAmm9QP5U99szoZ9WpLmURI1jvNZoHqarMtXsGMk0pNRyl
1cqOnJDppIvh5FW0JhIfXI19vSzrsoHHLGmHPbaB6HUtMdhAu4LB8gV6CFNVq2fhAl3deoFQuZSw
KStw/ca2moqfMU5AFIaz9nC8VK6TvJRZY0xBRT/+Obay4EWDPY/8GDAHeSNuQ/C1OTApqizdQAiz
DmhbrnAxU347n/W3ZdYL21ZXOkuV/lIrcX4qPg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2960)
jL7FMN9RTOQGIIN1qVb3YrH2p96EExrRJKe4eqER7XGR83PcNKamOUoE6r6Ts/+xkAOWs+UEtG5X
Lszfk4uDA67B/tW7OT3v/POlB1jS8IbgM9Hgqrn35GuvCUwqsXW6boVR5m4p0ZjchsgjpUIY4T9b
Fwpz2Uh3VWm+XQW8Ma2z0enReLVKIBnrEVB7X44Dp4X/EPzYDxd3zGPA+LgpJvJJutqgxsQmhQQa
qnp55GdawQEBBoXRKZmxmfmVPDCim5pbqLC/ZL36zqRNrzDZu2mwMFhqPTJ90kI1Y02K7HvDRYcE
gbsGBmI9oESuX3fdQT8W3P70TIMhbREFU/S/gAjPEu5AtovGbQCHx5w9h1farXLcsRl9V4gcqe8N
+OV6+4vTPR+grkV9MEJ6EWKiAZttS7GRS06wcg90VMHwJ1aHpCboC3cQyIeYdvjK6mRpKmQiYNcl
wlSPvzJlsN6iI1xl34ftRtsBVV4JpuLoS8YdXnQ0tqOtYPk8UW4VqAwpo4jUXqPLOXgAbdMF34O5
faulH/69amS4YoqQ9zWWQAiha/a8CXW76JMbZG+sQ8wNclqwq3IaEe/lwKt6i8OLHVl3MJrVFHV6
a9IXehJRwhf5kKOFrVPIYA/tmMCfE6wYzyL3OsEzzoh+oLUZW59V0qy+sxb3Wrzq4wpSTxKg0eTj
f5TfQNsxQI/guczq7Q/8yJ5u9GmWA/dkqDIKuo64JFmQmyUKIt6HuZnYLlcHz0qWaI5nmQmLOooD
0J+fmck9ZeoDqV30cmVPLSH9NE3RiYwPB0ifpwPQ4esBh1J53KaczvU1NbMACPXQmEnb9KaCCDPd
6FY3VBsiZ3dVE13dy2189jbW9u9rudU0L1Qa81qxnHFhoJpWbRmlzamx8DQ9TOYpZKpRiPYsMGuY
DcC/O1fSaLJFEFZROnVtW5T04gMqkIgKqY3OgNkuiyi3LufL3PlBdk7wchnHBodjUbgYry290sS/
SOT/zZ7TiQ9zg3+PfLdf2EDp8YEa+hBNMh/st40/a+pEiF5YlpJJq2OKz1yKYiAR6/ooj4/+PSc2
PI89iFwPXzitQYfCrpu/GH9nMZhPulQSEgZ6cvsMrv5OpX5j1pY8i4CE3IDqGE3kqjx62TlTA/bX
Q08LImHieQhNyyrrWrhiKtpbumhlzdtGbP0lmQ9lpvibjcR175tWyVmsdGYqBmD7HoQADMwY+Iqy
BWofF08JrNJJoTYfYie31a13igURCvrWm1DEuq1gFHM2WtTHSm374Yq4q0CNfex4Eu5X9AzfDDws
k6pyNy2jLTixw5WqmTj2XvgMrL+P4NKonm7Ix2sjgABeTyF6fGvQy68EIhWpB8ixprYCI2aoWXRk
X0E6IFgK/FKc3pgeTCo6dRGuojDRG5j5m2eS2WlCIjI6NUW546bLND4isVUU2LrYmafbNkM7+SmH
qglsbe7tYsxPUsAeWE3ZPTfWFASjzYF/65ZugBOtELzhGswhGgEYDB3nUQZYUFK/1HGuYbWxLHVK
wpE62G8IOMT8gbp1RvfqPuNCkrlsVq14TFFq9JrkleKOmri13ByFCjPO9VtWNRw7aY6aOEvJsVkb
sIOdEBEupszP8CQtJk9qsQ93sKrpifvRWBmfnAM3tvFppmo4CdYPPoH+07IutEmgLmhNCfnu197T
MS6PnEA7mh6vIK3+XbOFXpsPA4H4cuMR/OH3qpF+MSQpa77VYsA6Re5SOqQh3rA9XxMfy35Mynxd
c3So9t2h6pa+OLp/MIrq1MfvDyxF2u/F4r2Zp7s3NEElZdj58PypI+I7UHofllH0IyezbiLci4Oe
x7wkYRulpUt9aCHGjw4hrWKAbrm/r65s3hzpW2Qseie5txeERHLPcp5/CgGP9YFZCtIlX7BK+uF+
l9VDVBafl+/ZxlGlQ6TOmjf9zxLOGksOI+4HAVjTwJJy+93G1MIsq5JOW7gg8SOMX06MVpDaWfmZ
Pfqt5B2wJYogIig3XAdlpe9mYqLZqkkwI8+rp9ylhxyenkNClmYn1QvwJ1a16nsgxvNKDVvJ83NM
2+zCj5r+O9Lk5DmCehA+y/jTzwvwtkHUrE7KHxDVJefRtX/mp6EiyO02we1ZBn4+BtcwQEIUrCBK
l3e0r6+ml1WXmUjNwBb4yZ/uwZDBIERi6csSbRhQMnZDprSJVi28TkMGN1u7+x7gyHjhVSEYxM9d
rW9DhKGZXE8oiL87pirKQKWmlc7wL1WOyDcsRoRaPKYz4K3ltHCppWH8tnwbxZrAf4qDt/rCK5gI
B5E7go3zXwxLAYC3U7oBSCrG+WLY94a3O7g3zKDH1mS8dxfhqaPhBmMpmVB+DgKDbECNyYEk0ddy
CG4yPuGNWyVGKEm0tALpRFzBiCiKxV3neLNhJD6yXm+CQHim7Ch1Tjvi2kM4F9JiV2mvt/+jAQiU
VRXW64mH412fkqsMQLv5+BhTE/USCL/xsUDa/lqVbX0pvYyYsn0bjqCkWPU7Hg+Xdqj29HnwQYI2
7OBb0bnjzWPmzW2pVSt995qA2a9+0AWE0cgXHtGEAFuOqfMg7JVfvZmXlqbeKXgyUCNcZN0xUsKn
gxwIUxJampvDGYGO9xUu75XzocJOyh0Nghs1I8ogOpixWqV+917ptvB+CxDaolJ7x49YHVEMC9Nd
6bmBcexfaRzEDP6GEmFxN+RPpqNr12vh+wF31BbpL7x48gg3ZSSYRHk2NaN84LxRKvYVbibJgIUn
hnudLFioXos1XHNKJbqL8t1Z5WzbSh1XyuRReym5e31nQ3HU0GJv3mNnfwyK7ms4ZB7JmFMCYC3E
49BFadntYEtegfkkwKocRwvnn63Mi9PQDyD1aKU8GlWMrVln9a22D65aHbzNE5zGw8KKrwxoB/Dv
92kY2bWb0OiPgPLkKYCTrR45ObA69OYjWb7aiOu2KdzFN+HeIZBNUVVDjStO3VwGXtdeiT1qWq6w
IjAp33lwaznki4hSjXrjn2CeE8uk48R3mh7MmttWZObLkazisPzBj+eJZHlVMv3aHZgI1Tc654BF
hU08+7SdRCgjliVHppCXFnMxFZDiJw19MDOL02OzpNE9rxxTfcTXkguCd8S+trazcvcX2+UCn61p
SphQsyLpohQMtYcKY2FanqSsfiLYcTyYvHVSIPcAgEAcmSSSQHkImeRBE6rLQVORbslEmCu+YUlz
NGmpQ5lVxRrEKJdfwpsL9tVzki8H26YHaj9yIY7odCbA+hIx4kiKJoQnlk7b76/tkBikF4YnNrg6
Az0ILbyyG2bO4OAVwyC71EZIgd0JHfueaz4zCCwglO25kayaQl6AQsXq8r9NOKkLyksN2X2H7C9j
5uYaepn6vZ/ADb08nnie74NIItwNK0d0c5fmLAu0rx0fO8gGyPLPJVGAd+ab/zp/GYByIUSQUUiR
TcXI2A+SfMT2sseq5l0485lH7ljpnpsX7KJrhudX6U8m9I84mj6ZMuyIdKoype+PbrhEwEErfq+H
9zRH2gWshXxdWlsWFnCtYK2upJRe9szC1CO2U7ADpLR9di41cQN/W7FLOwUggdVSv7DpfAIkJ8Ql
rSTJqbgVTDMQ+fpdYVjhMe42hjGJRW1/k7Oqm12IrudCiJTtNIgc+roLt4jp5CHjDSJwcGX2CGiM
ZUNip7b/uGdN7l/a8Sm3qMN+//P3FypkhUp6XB1FIaDYjZNojH545WPdekSaZaLgmj9bxRSXhdMM
rLUr7dzkVdoZStBk0QUuDfT7khP6FDHaOOrA1cSV++zLDGPkIPkIQcUkJs16Lq9d2Wxg7US0HgI8
LIFyhjoKpuABxSHPWYerFeEQn8i6Pk3Bf0xVdrjjTnhQpQqNdj7egHxI/Eng+JbI6C+k2mgHEEs+
w+BpZq7o+DCLYaJ7jdoiSWBT8WmBtKsrOqhXbG6k6sbz58f1RF7MYEOkHUiodGvZ8Dbm52w=
`pragma protect end_protected
