��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��y�1��pP'�ϟ[�{�u�su����.#ĸ���}��e�C�jܩs�TPb M��kw�0 ���ztCΘ�q
jO=Z��$��1b<1��3�s�^������88��q�r�bc�I<�L3��/@�����[IWdY���Mj� 5}e��"=C�ϕ�	�?��:w����1b�OPsdT{���%�T�q��c�\OJ��:"&t����w�&-��J5�lE?��!�E�F�5ݦ�؎b�t
'���5B?B6"��w�r�E�� ;~�����h����.�67����$�z������N/.��� <�̹�d��ܚ�2A��;re�p�=(���ǋ�� B�Y�ht֧�*1���"6�y������-�	�Tk�l
���ɲ[�Q�8�
I��]��
��H����|1�G��ܦ�RE�i{��������^��gW�'3��ƀc�7?{'�ë���P7_#م��jC~�Ajo�Wã5�7�wtb"�Y�HQ��Ϊ�C�Y���?3�����	��-V�aPr��R�S-�=	��.h�U��|�|�h�ԃi`����Ћ���W+4&
c�ݳpA�xh[�I���%%������a���`�=��X�m���C-p��
Y���`H`D�ƞ����w��|M4@��1�V�-���(0D�QD""���
E�ML��3�"��ܸ���	Ү"4�\eQ��%#��~o�lzlP2�D���6M���X���Y���)"焦6E����L��q�OE�Υ��K��W /�<��m@`�2�"��OrM]{ɋ���C���o�p�>���e���� ��0+����0!�C�J�뎪aS��s����}Ĕ�b���E�X�(�\.�t�(C����иM��1����c(4��/��(�ߑ�`ڻ$�}�e��t����J�>�}x�b�~�����.��C�:H �o
�G?�?��.�:�~R����>xY#~�q�?R0\W���G$c�ت+�["�v���� �-'�����,�g���nra��5>�a�����Xu:��)[+K��jH3FB��Z�\I�z:n���n
x& �Ww]LxA/{ZR���5���U�"0R_��7��;�%f�T���e�X@fQ�}A���6YО~Y^̦�dA�Փ��K��؛�D�H8���u]|�x8M��2�T�{�%����&5�0L��H�Ȓ@wĶ����q1��Qq�G`��H�^/Q}��<R?1��0���?S��8`9\��H�����Ͳ�sK��8O�=��vz}х�Z��V��x�=͒���u�7֌�#�U��^�]�5{���!�G���_^��=�ˡ�֌�����tn�� nT������`�5��bBHXy��Z�0u[O�����r��Cݑ���	���u��4�mݙ!�̷Iej	��[Oxcnk�H�y���#E�f��I����#\��L�i��.�'Q�����:��+� ��.f��˪���� #�^�@}��LO�w��