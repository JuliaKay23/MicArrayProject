// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:15 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JG/QRBfK0q/fImFtPnWs/Psku0D4K1Wc3JPnG4UnBOSEmzaCAaDKLF3XUNMa/aBE
Qman3Wya6lzo/JpCU1ic33/cALCMdTFpw+oDrr+GbQUAC/Hds2YoEQSPrRMky5QS
TQbxI81J1bBEkrNwbs10+juO0/IHRgB5TQhKL4kvKbI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14080)
f8cMwULuOBxOPr6BrBBwIdMmYlY1f5WC9F2pT4K+7Lwv3MSn+Kw4U9BcG/E38FLn
CDAfCfbTWKRb18KcUjF1eSrriU07P/zUlqwA17MASlBnaebSA5ZB5ZwxZhrI220f
8mBUjdVrOWLlxB8TWIMYvwr1fWq1+hnY9FhTLWT8wZBdJNnprR5rELCNbFe1dMIn
XllxmyAz8wD+tF71D0Sjne2nVZcKT9WGQ3xEarQK0dzmU81S3pVTvJbVZMptpxqN
f67pLPYz9os8fdA0x3DLCkjpZvdsJSrN5jNdOcIpickHCHAtblWfvJNJwv8X21k8
Cf+vjPuA5Z1QXMq1/u7WxyZ21+WNao9ztPiX+ngZDhJOELfLUCjNPBXworLzTBuW
yDX5vE/XcRSFvtQVeKJPyz5ZFFpYAeOd1eKJiyAcMI0NRnFxMnUJwZRyOpFSr6TQ
NwX5WYetZMxqhkUzmrSZtxBCSsFLX3U11RFueYY6mP5GCEmFi8aYsqQ3kWOzsYHV
BaE+LX02eB1kY5949HJhbYH+e3auwTBiw7LVZaC6w0nvd5q/D5+y9PeKFzpJ395p
42NJ4LHAx64z6NVoS8fw+uksqjIar3MCmz0B5VubmHhSBfu+pbegDv/k4RvGxJZC
IHABsM9k0eZqfnw80q+kGOMMZgbtKQMgT1HPBZt1VVDnaSueLlniIX88YrW7wfHd
oKBzgJhf6MGHXoKAL4ufsg9vESh9y2n+F4xQXfv4v8D4qy3CbdeBScRISVfavHBG
aDn0Rp7crB5xOFJDXhHDvZsQYjWZLk+7GczLb19PB589WO11WjskdsU3ZWQW6oA2
hH1yfzpmxR7JGqv3fEx9reBCYKF/QRuv4HogoUpkQNgX9dBqHljdugWE+DbZZsIn
RTCz+EDwZEJOAU0khtV6W3ilT7LWTLAMjOwjK7Jh7V2DCx/WeDvfJs8h/MKMjyOg
oABmEgfdepX7j2NFExi/7YyxtTHd2N/vKtfd/fXjy8XLq8eIg90w17XeULsr83Zr
vS/6RlgxR1zK7Bt1H9erMqlbV8xJAI5TyFVj9RGabo0f7vcgJEazEZLIE5ZbwRiA
471InzojafCT3/2VQZ9NbqzIiHki4hLzoyI/LzooOqJSf9pFgUmfCXq93ZCKrVqC
/fIUZzf8S0VOM6AXxUP7Ge40o/Alt9SzSD5EKfO2Y+H/S+ADGHkKOCT+6T+S6Hud
yDceEUTJcwT4Rr44VnxPnAx0zaL9eJ7I5qDGoP2g6QxFM8+JkqSAebSZxwx0CS1z
SBBRTtVZaVvw4Ikb3wORnagGEl93qrJT+p13UptIa82Gv7Vvl7U7FsC/lpmjrCMM
lDAAhn994CI0DAwe69Tz6fOTPWjtGdBbMYuLZTA3DKcUrAvLqOxh3rcQoqSxZC11
y5E32Jkl7JEGJ2f25Dwr5f3O65v38OWw85Qmbs1B/MD+eDZdILsmuFYsWwV2OZlU
rSFOf7kP6sL3/3Eyqhc0V+xoaOt4Z+F2mob2uyLXTu09IEtw+DcC84zkhOD8vwAx
XrlniNOa1FP5vDInbvZz+iO9wm6c4UntN2dFa+PEURJPFrUmI9VNBrJXg9quQFX+
Ork8psvBK8Dp2t0haVD+vkzZhz1fNeNNMeFFG+IqmzZKs2mFeH8RspqCJ7wNPhQp
uvXrT0Ffv0IoVgl9LBvAHx5pi7vfDyfkRxztp2OJQfU4s3/IItKYjux/ZI8kOrDc
HW8bnj8XGc49VWBd3+Vl6m9TlWGrTZJVZ4G8rqa2uLkBxeqKbKKvhD/dK6550JHx
D3vplhG1AhnES2rDLezRWhEverj3gz8GN14E6q9GU47R5KQlKwMIgg5Ouf2xof0X
1OSh310Af8CBWKhv5Th3Cgm1FI0Q90b/HjDpqTm0tV0fJUuJJWVYO95XY7plTy//
thVmYjhL0A7V+gIbikuwlBBFQODAad/kUoEYNoFmpPSHxbSdwrG3pOWh92VBrgm8
sYSBlblUANfHe+AnMciQs52TiizuOPDtn/bdZJEnK9wwR/i/Dqt8+Kz69kN+JUEd
83s0A+886QxP/TpWspk7EHNSi8Nr5pmXAgBF+SkuFcILFFLyQ944if35VVe2oCv5
7XM6H/Mqzm3YrLgbiwV4dNFy/d/KJUtp5RXIa9T0++E6dZYjZY1dbR18zt6bEAZY
Tv64cYs+A5vYsEqofc3u73aClTDvgmh+dM5dFZ6ttCLkIWZUTvU1ZJPm8w1fEzv6
OJW4jzS6NJbsrCbcsOOIeu2C0Hf4Nr957FTgkR6pSkWg9/ga/oM6gTPhShZQ47Cn
CvtEQmr65YEMCVlk6J82/0TfQPPRcT7Wn/FI3DxoY9HCdtCjBiE2tmq3ycFUSodl
sOoxI3DWSf6muDOfqrA8b7qpPoIAgMGD8qehKIcXMNHX4P2RrcVWTepLGmfKwZd0
aoqzdJhaF9NzpI1U5i4JeeGQ7MJK5S6/3P/mtYnRrQfPSi8QkjCtPpd4OpePqSpt
yQ6uILLJ/8lAYnwg0+cl/mIIrO/Zh9XdJfb37S+/QX0GtpiQDkDEyueJyzO167Tt
ZcdtSrS1v2MvJYpkZegQeOR2IkTDsJWyEpdHggs/X71j/vDM7ANLtba7z30DQ1Ag
sS/9dX+OUgD6RpUg/VlAzWJXYqLTBWCANiXi5SWVeU35tHhj1XtcIl8idp3NmxJ4
UB5SBdqL7R6DxPDMhx8j1SGwDtB93ExQVm8DIyROMOCld12vQGokQ48cYfANgTOE
UXw/0SFv9qMXPumwCDk0ZWXAr/+S8ZPy4ngCwl2udQcHWiZ43+CISaWGOglLfSBf
cxeDJuIAnjuVCueMClICtYjHKiBNRUDvEgDDvfzWyE9w0RUGdlQnpfEuy5MvqlmJ
BFkBiD/Io0dI69ZHKyxQ4a1lkxVTV8sdurqJjz6sCG3AhO/U618cLNxC8cpqCc+k
UZXCnpdMAQDpQIDCGrhVmT0eLePFRt+GcLauuWxVIKSxiyjsU8yB4SUI5ffKiDtq
qWVpKY3kACOzNYLljChxAOupx54nuUhTDK4Zr2YgWeBOFetTiI6xoJxEk3IueWrn
IwMKbKT4cgQQe18kWC6e+Vd73nYkgptglP+S4qYowg8FeNJgTIplYR08u6BIGo3v
MreTMbiYtzi27aIuLYHrI0J9ozUvHVUnHOP+eP2SbVVNpkzY2ZxpWqxukwEzmDeo
kebn+6TeO/z9JuGRSVDPy49GsSOa2W1BfFT5gjl4CUvT5Ny3U0aI+PpDrFnmZELA
CD1ztdQNrKrPMpGbYwPmXjtw7u3CKgRLMiddDxaqgGOYTLL6QudP6838ThEoTHFO
b4Dv42Z8bxu/2al+n7HAp4gQbS75S7ANQpjW94HNZ7p3MecQnmq5vDpdvdVzTJe3
Z+/YOZ5VsDAia2JOqJGi2BVqCRzrF/fweDO0mepwD8B4o8LHwNAyu4wF4HDcqpi9
05FOps3gIwMFOWxFNybdfYMwIOJXhO53cD2YJKZd+sghCtkzTtK1OWKwKNhnH5TO
QdOtW1AsQOS0OelvWPB0+5mDz5OJmYmIHKzTM95uESdsY/ULnzfoKGlxHYfwWtxw
IP4356EBrGigKYBtGZIQMhriCcDGrqG8JnESa5DPCgihzn6iGjzu+YHsTxy42SK2
fJdl6uTviXVAGt80S2w/DbX4a0oX98wTBsuT8mpY0h3VNr3yoR1BvWhIwhT3CF/p
94eN/lkqa+TkLn7gs0CdYatDPxqecaXMvvXiigfGnfd9xlebwDWfMV4sKATmnuZl
LcOUuFC5vtXT+fHs3H0v3NLPyXlwlakqs1kWf8OOqKa4djRrzubboK5a4emvkmcO
E7qOgdttcWKqRGVEE++7ROf5YJV37MSZ+sG2IGbW3WQg9oH2umvVWH/gO1+b3Q/x
ZEPudPOSpaV/eIwgTG5zG+U6CZJMXChXu5oP+88f++qRrM5nZ2WSSxC6LPl1genM
z8kdpp/Fj9sDZ2T+s+EOOMIgb6F9l7VxHQP1dXZQGeV5qzZaIjYTmgBlRi5ENJ00
n7s7G87DN+3iUPE7T2beQrzIFR5xHsAUIAeV3t5xU5uthbbc87zGgEPSfpTL1AsE
UA2wn1K1SDw4saR1IaVW6Z4Mk9FgCvavsUE6wQs2Sb6mlU+at3x2mEjKa+09QBL9
N5wHVqelXPldN6FAmY4xQL1tHLwuyhv3E3NX+KxREFwzjegPVHzdXZ9MlBeBtXrc
7syRZgUH35WjY5/XsgB7Rmy1vhVt8brIeKABezJERW8APySMSKJkxzYhTz4m9TRB
fHSan3EJZbDfNQ9SsctxN5qFMG5kcE8rkCeCcpP6JuJNiaE2pR/bauyb6mg7718M
lDqVVLX93DEzLW+RQMVD0HzcnULAeGgYFfBhaOD3D76L1pPpp7QHEfmlSp0APifP
dGczZd0wVHKQ8ycm2MaQNEOQEj3tuzPjGflCwxhns1XhhabavyRoe3TDxVpc8Dlz
Rqlb1rivDIdbpWxytW/v6i69176VjzXQ6B6Fu+4xkUG6mnkM4rZf6OQSWqHV9EkI
C/k4rIRbbT3XjQxdexd2fZiXhwJnrbSSYSDYphZ+xnfmLv82C/Wnv3LJb4AzrKmB
f2aZiQih4S2v+kYLMyX/BXU/hDYT1T1XRcPwGyoLJRczWJXxOiYyRMoZVUft6CFs
5T9IpwfS4jjUS250mcd8uZslhRIz/9w4XYwz0nxo2iosMF1UhGkt+DV1jUoU4WJ1
Fx6AMQR9TyNJCouefruit1NpI2i1mf2AGrmUNWTRfX5WNm2lx8mv5JIvwD622G9A
8ZROF1xKnYrIDFT1+scUDnhGDDBI6ulW9Umc1iuG3meV/9DJnPo0Yg4XxzTRwIiO
265wJwFgwnit+VpI+FJEiGPGvXipnnlIT09bMfnsqZXHyEGek0mh0DG0iDk/gb5z
+6wHFRFZjC4KpTshOW49XbP+X615jk4CqxSZQYHgfF3WxvTCgVdXQjeHx+hnyuhj
puARP9ccXzqL895VwfXt7pho/oq3xlHaETwKR6p0cRyB5giPEOYyU+D5unn9autQ
NYfbI+sMEkXcSkTYTvvKZIFOsgOQuyTP+jWqjxSrO22heum2eqmfzkx/X3om+KcL
vRNIzjD4OFlOap5I+ImF2/3uds7cYioRzecycU6+s+MJaJ+CFIKCtZKKIoyVgF40
7xFwGU+QsEswRDKQGgTseWjgBdzGE5C+CcNKb7beuBaQJfKX1pKlKSobTXT/k5ZG
L6F4c4S3Y/jjMOJxotgA213ldcEO5NUiPicLWyf9/Zeq9K/pFJb/pTNb9Kqmwa6i
FcurhCRBdys+hSrb8RTXo8OljfASZ4Q4FEp8+q+YEGOWdMIPA2JzdgJZcCpAzMqG
xGKJhjNDQbNnpLmHxX3n2dH2Y5PDsRFIQD09OofMp3JpR2DH21r6IX0ezHLStkKT
sZudLg39WKfJTkRHu3G+1lHDcpbXoddu2uQmGoClBlxPlCM/ZsptSbSOr5QjHPtE
2Sei3bQpl890ZoJBFA2vpzjYlZQtGl8QvWBpbLNGu3XNKCqrv+URqy8QM86qBSC1
EG3VU9nynA7+8HZpQQmnj9sv0zgLQRzaV5oBL+M3w9h85qUOJ4Jr+sBYojoqOZX8
E9Ia0ana9h4Gg4T4IDh5EzlvcBPy4t5OcjJSMJLUsRkKXm92C616w2Bi2njmJ+vm
f789EL7SUm6wIEUQlnbVp54bQysm7Q9GTGLrJ8LhIbJ6k0UZVpnus+TIZQXiTQDa
pg+ECsxQk56AQ4V5zoc8WHv552M4G66Et0dD8VU6E99c+KuACX6LzVOEOFheKuJb
oRAFA0Fdt/rpW5EYgGir98rZmbrNlQxn9YGCK/0i65BrKH9oVEsB6MBCBwIxbHO/
etDf3MYUnfqq8wjV+MQh1jTd4yscQ/p2lM+OZaCAQVqKzuItyWQAYOPO5MvisWiY
1Co5W/1ZwHggJEHwkBlYd0K3oFZh+OLLkcWA6CEq/X7FcqES9cFSSgZHlDjujOxh
8J+XCxDdy/LWV2Jc8hODh6JOP/kpOwjEk/hbHV4lmc1ThrG78PigNxA8wv19DCD7
j3qYWuY030tZwEUgGfo/7zzL9ub4+9gXsRsSX+LG0CoPOUicmKWjE2eNodOmfe/j
l5fconh/AJLeoM9DnMgnZYgBTIdmk+TPlZaP45w+a7Vvlyk14kR4xGlL4smUQZXX
R/E8u+i3VJzBAg1Q9S2vnrglYl0tO+UUVxKt+MD/pkJcw5aLv/0WlGgA+1k4XYj3
JsKBFxLFMap4+T1RNkq5Yr9JMKEpwD0Q/ydaqCytNI4erCKQf7dnghuXMPbfTISW
FIZ23OqEPPSCk0cfQUobA7BWI+Mgk4c0hWKol4KIMCP14N2SaP/uI5vbVVirqQ1O
z2Tmb9VNhcisghhTkpGicUchWgXBHeicUq451Jztv1c4SxxBdBV5WqvWyiVEPjoY
oTz4CrnJ5tld02LK8y31f0xUet0v5OHwe0W9SRawNN2o7naE8jTLCr/P+MPLan2p
AQt23iYByhdBCfBc3q+uqe6CUlsV+R1c5yf63lK7IZZu3IawX+LF1hwDg+DIPriN
Zs6TotuES7O/RYR+dKTAAI2CqnecMS9NcGuTFcS/ZiB0v6Ky+zIBDySBTRjZafXJ
K8LW+cM3CX7KkVj589CPwQK8BIOeKBUM3KAVn1koxUWjIYd0B84hhJMsXLmUBrHL
v6zreyDz/3+m9ekQSx9Py1HPPjf+5cgHGOqxAypWsL5Cvf/eP1Zvj/ivflawCrQB
JjDhDz2S2TSZztg7DAonz/5gnvgvCHHD6kGwitavpMjQEBB8wyVF2h3VOzlvQBpv
3GK4WfjsrI+VHJj7a2+tSi0KGKsAUkiLEoG6CWpa/Ok6FvP4F0/AH4BB92q1i/o5
m20mDkGdZYkMWjJoAVM+VjYMjhKK2fC2JrlYX9B2WH9rtq9wonFqA8E4jErHshLJ
0jbzXjrektKLFx7SW5PoYZT1w5z5pYAzmn7J1yGhx3dTtiIJJjQl4l0/X8+qVyvH
0DDbF0Z1fNLZx2gGcX5piGUB+47MUCMr7/1vCXD0ynm+47OYTF/fYIBTdhTrZej8
u6PUz/Sp3Xz2DZscZ1eAnyXGqCXXpCQTHThOSjUeMPJFX/prxKRZx5nUMPSyaq3W
KTkV15Ec1xj0c44sk9KlX3TfcGPy7J6JouGaUTfZtiIraAAGZ0PCjpzkVJPon7XL
On2BDDoiCdFelgPJns85NXb56lzuqlJQzt6bYfeVERl8MtdiNwY+4ti8JBtsLt5s
mjKPlMV1Knd/vzmOwdbNE0J8bqOT04A+H8//YubxqJdYimbynw5xgLfznNMT/jvG
wj+CsZ90XuRUYH3vTFGx6Y9jI0PNVCq0MMX1Z9bmCICSPHXgiGri8W5iW1NgvVtA
v49ys1DCzweMbCJBLFEoKbL/rXrysqpIK2qPrUG6FSmravZ0XBSMtMbEUmeEK9zp
YOiPxtROwhv0OfmHHtp35oIbhVkZPfwzaIDbCzjqaF+nOILSreppntCcTwoh2J/h
XenBKWbtuZQzjEkK+waKR2x7Y0RFp+TJCIdaUOwVlqOOXsm31xvo75BkjYdrGNm6
dv9C7RZUFAQrSxwOSUmHG5Du4qqibigIBo04hobM+zBU5Vs1F2qYr4RFKIGktoun
ItIqfeBP8nBYBJP9k0pWXz+L8j8PwS95LS7YJ4DA9YpTVkfK4N0ClnqHe8AETrQr
AVpr+U0DuDa9do8fd/IsHsBwta7rKlNzrx9P4XNaagpEQ2A/9pOlELHKxPnBn8tK
v6PHoPAVCgj29KW9y8z001jUWGnbKDYBCn3QHFiVNqrk9E1bUuFdKsTidWTde74m
mZGIe1bzMboYeGWX+bKAGOUvBWkGBLm4AaKFrq7nCJIAH/UkVszylDHARgMAKgTS
LmGWnSYdxyRM90lgExxjo2Oo+GIasH/WkWhHQc/UvpA+RSerS6noI5rpZ+a13R+q
eIiBU4Hhiebq2o1W5PJDfIZhmAtLgeETDzZyG7hCGiqcbnYRruz42AflXOAmYfIq
EJO4tjIYXBFGWkei6ht5wvKsYSm0NoOkvVOblDfwK4aRigovhI4nN8ssuMSie3ro
XCprQ6AosOOsMc9LfAyK/3pbb312Q/jRH0aMarfAvo85NXH8fvsAMpaYr20zPv9M
aFX8c5i4HJXPcN7Xit7G4dTG+PQiOlZBJBy1/7ySwUJz3NdUyu8cmxkQG84YYoqq
8kwYx+rlK1ybQ/YSySIwmrcpdXK0T4rrtdCc9VL8+m6IKCIkKW7VDIIhWSOwSCBm
DNeDSCS7fbibjBi9dGDt/qW/cqTmDWQuRfiYii/pGgDnURvvvXlnLYKvdHC/3xn9
nULetlH4bc8L6JR8g0OKcv0ydQkGVBF7X6oUhYGMf6f7/RhrydEaXC7qjcIt7BsV
oo8uVZVUfNeDG8B59cw5LbQJAVr4MNm8cKca8xMX1YUiJdrcrJ3+AM1vDDPSzhlP
PpVDZ4ZNwsvLK7K3QOnFNfCmJkfAvsSe6rKAqdBjSQhL8hN0aQS+ZOHTL25st53l
NMSjf51KQhTGv2sd1uP4XhxGzlbaRkoLkxs1EhfBwt/iuAF3aYKDZGfxaotiP4hD
q6dDO8e5hBaaR2y47holSAgFho62zSVN/4VG7UcK8e5un4ICfrHK6xFtYVq51hq5
D295xfkRdBT4gZ7MIPyCPjAXMLROKKA3Ex68IDMHeB6wLmADKvtVd/LSBSf4sw66
JpwkZthLAH5SKdb8p228Ko/WGuRQcMQ2iKfHhGXoFUZADArwwi4QemiJYGYAB8u8
BdgPGwv9wHeFajkwHpxUMpOb/3RoRzdhPYuq97DeGzCCpFWaoIdbeFN/zaKnot1T
YSaXfONSSF+IlUcOEEqFBfrYw0tQ/FBu6OUGzg0wVVJmKbn3YzsQySMg9rQlJcIQ
bMzGYrEwUXdNp94kfJ0kXgfCjmULDfMdy3C/VCgLc5IO+xr3XJOEPBi66UQDn0MG
8rz98rAMun5sriWsqLaLIpXiQi4S0Yeob3Z85adAjn86bcf8N9N4o/w0/XJi5jPN
z0N8KIo1G9jvMfaNdnCV3oJ9+Db0/cdUBTGY4W9F2CauEK7RDFcSX3qUk2TfNjee
xVsjaWyXcehG7DEPCWU5LqFXO8g0wK5krxK3Q19bF6h+tPRVrBpqynCXSXsnTcUe
/24hCj2vNWL6ukjoykydw6yYcHGMydBfmEQsWiraWIK6S9u4dAoWvZ2mZgmeJHKz
UbA4UpLgkI95X/U8V6u2bY2ZLtLNf5xLx7xbaq92FR8vJBuOaI888+l1Se6S+W5J
q7tjWWz8dNsrzP1ghh2oENIOQ+CWdjUaS9g6XvBkk7cE0H2kPX15C9F4TN9aDsCs
pjLWWmrHd1nFBvjCc+PamY8jYVz31DRdFI+x9LUCqw+gbhcz2E3O+oW5DGrHxLNw
X1Ab3pEmRRGrInL5m9Hx/X9bfh4vyx47P3nZhnENwqj/+KYZzsBowfFgT25kI/aN
M/OpJrdhhOhRwKOzVT9zr5wO2Tj4FEoP7ZkNdI/+455T6A4XAq3IgMMXVsG589PX
uQ4rU5EKyXefUzJEVv7Lv7pef/e3+Y23qlbdkque7Zccyu3G1Uz35FttqRbx9gH/
aGIBIoWvmkUngSFuokZc7ak/rrgVqn/or1v0QoCksms3QhnGLGINDxn189W8iaDO
wa4OXmz96RR6L0H3qwbcZaPbi+NMnNLdE7MuWbd1ZX+2TdUe0O4QwIg69/RZ8TXI
2NkDZ5xqElqYCi00i+sahDebyWwgx2mt4fi3SvUAK6FbcDPVSDiXHgGvUyPlc6xs
KQWiWqMqKXoQ/CuWUpgM0gqighkQabNi1Ue5Bf+aULe+dEnefNgxc6DGX2SpPdfl
h77LVbCqSAEBMwj6AqZyZJLqafwCn730y3GfIl39kdym9biyMScLI9eBAN2aegP0
rpiU5mOuw1ivqKoOAq5k0rJqNclJX6LMYgjGOkTScWXwYgqXjiRp/lZiTGj+r3RJ
JVEz7RfuMCbKlQJMiFdzxNMnM56Xz9QgRBHCPewGVrHvYpSSIywNdCGZWLi+eg1w
NXBdc4JUGxwBobJ0uA4jvTuTemx1BgGMaLKn7WzhjNqYA3mcfBEqklBl0tnpUveu
32P0qgSNT1BK34UKNrB8zT65r2pdRMOdPxcdO0+KxWxREFwk62geT5mgJKuTGtDx
OG3G+VabNwqFJQe+fJXOGdWmCVuG0/8R0fX36kGQZnewwvQhl91zyeeAGPUfLC3k
tRAcDD+ty2xqCACEmiE/Rwj1x0fnPoAi5GQxbp28rMtCsAQnIN6Na4OleIhKj8bU
WmNDAjXW6TJ30jVHWlAl1LGrSdCkWuRb/YIWf7qyowEsi/9eAXU0CefxFGufQDLY
56tIw4Clwswr2mSFB4NOPD1DYQAEDlYpYBsx32ADTWT6L9xNnLQLfC+ojaNOsgGp
fynPBl2PRvJFcfFfarNhP2c4WU1eyudmLB29IayQ2FBVHv0R+cDMor4LKP0NcV/O
XYc1EzB5F/5GUShZofb+Z04LMV2YQd+ZLZGg5JyO6niZuXoFRKp1c4tRl9wi3SAW
Hb9lIZSE5E3nTAKnOoi9+UiRDaNbk3QhdiV+RlI1Fr2pV+up2xfTLUKXbcLIu8eS
hLLEaZjsEhL2XKQ+piUybJsTt5GzDC3w4LqAdKcjLhLejQmHA9Zc9fzp0wO8XNbQ
89d0FseW6xwEmNdeZ+0qlaCMkxFygt7bzLFni7QSjX2xz7Gchv6HasavKv/P+x9f
XFNOG4+dHeRuhaIUraInoL488HTfXg9uav3HFjGbisbvTfrDMWEjfL9ChmY7x0tJ
J6sbhqtemGwkq0dnHd6Bek/Mv9GfKNtcX+ILo2dXxqP1bPRVr1XyUOpafE8PpBkP
kx68V3Aj1jrofOTxpdGT8CwhuOmzwDBA7fPbwvQYFtPHZdOUEfds6JcirH6kSeXR
CfGlzi6tiqjLLb7O9ij0W4yPa45S2QJxne6pXeNCa284CeBjg7H78PLQTquk+CvA
Xx375j/wR78ElbEhMZXLrLqxJ2LZs0OzUrArJ/lEmPAP+pe1ppcWW7USase3HBYp
KucbvyXEP/wLpsk0DPkcNV13d3KU4xbe+8rEhkhu/PbX5RnWnEo+pumT6E2GF09d
4yI586g980U/ZTKuBau4WQ1x7OdEFSLj2qs+MhEL2zbC77j/exuXEj46LnmfDrzg
S8YGgkpltnTDoZR03KtSWjeV3gTHnDHZEkX6FSqWqJpWNjtfjikhHCh82HWWH/Uh
vFPKWYl9jwwSoE2PctnNTgNgkqicrpAsKr9fNNOP3YOiT/58O4GdmlRS1GZdCUXB
BhfBvpDvMWXemMhGgDIuPnEmhNutgsOGKft/O/0fxwS/3CiXtZpF9ROMjmaeZ4Zp
k4upw8VcB/MMbFAQeF7cVnnZNOLceTjVx5IORSRrFIsYhYTbzVolDvYJjQBShvUl
egDOZBwFTYGv7Zj6+k9eBG9y/Ct7l9u9jQ5zuZVgCW8T2cFyf0r4raYGjXo6HInv
Wl/RZ7QwxHXSYUtev1QtRCNtVVkYI3U9vEUf6Jj9ZRtF6zjpdM6BCYkkZIqnziTE
64PGmVOgTdjDXwUYUJ1RM1t5zPqG/PmQtPz78AcrWBeelhg/RPuLZC8RXT0iwg1z
uCX8VrDwePEgJStPg2Nn07kjr2ZzqroajUSPXQ0U7QkGPrVpSRHj+89jY8TCuKvP
OppLPIKg+r/LRjqi7Ex6mz8jGirottvMt4GfO0gTg34iFfGEaWRrOo7kENJd/QNk
hdNlW8A50QF3ZOtBHuX9ZqHmKFf5nKKlyit5X5acd5psTvgSLIUGbJv21tuiUzdg
dnh6Fm9d4uuvNsElePAEToPqNJvR6ycVlsA9CtKrp4mlHA/PwlqX9wnKvQGeqlCE
6znoLn5DmzWj5oZL+Yb1llUZngCR21mACoTTiXhqlWncIGsa5I8bcsFtToSD2Idm
XHizXQqkbTeq0ZV+qbM1sKK8mNqWHosgkWRMoIeEgGPi542xRruWVyxxS6xBHz81
/5Y3WHGZidejjJwwbltkAZVvWPSlgpJvknUfH7hRWii4is+OP30492upMn6aWVQ+
4O6VWD1rm5lMyyrmvYgwc9t+l/ySE+PRC7ewViow4fCwOso+OVnMu+zKqiUY5Wo/
lLT/2g2bZ62uXEXaQ0SPYJNoB8wxxvRpswH4YNZ2oJMf8fy5yp0UZqbQq+4/Jtrd
pLpvBNpTofH2B1dFsRU/9WWgU4HzBsrKKrWHODbedie2oXCT6kGgiaiJX8t3shdq
2N6+vTLLBD5l7STLZ8qSHs5xGJc5PWkaUNz7j06h9EACDvYuoJGW4VuYbvEBNk5b
TST+WNGj4m9X4dNJEwR1dl7xgLynXlHKlBqex23A4Q1oy5xCzmgefmk8p9fIR7XN
gZ1ySqn1Eb6MfJZ6o43+j64DYmYhdBPxtMaXnGGOUn0LB+9Yiujb11DNc54yQdJe
ebqxVFSva2GTs3rH5uMQiP0LkeFmNw7iWKni9qVoFoo0YY5LvXlxWcyaa2byF1d5
/ULKSvIZw4rEx5Qv6+SWJo0cGKbkS+23yqvjfYesEZUhhdJEP1fBHKw2BgdenF5N
Qo6RMZVnYQr6ifjg8av4GQnD3UIG4IlJif9D+Ag+A0HV+QBy86mrlAjedn0dzdtY
McHsoSVhjoXsUf/8NHjNQ4xmgAGWFBFi9SKeGM+xtp32EzDPSbca4HfjY4rQymmZ
2RekTGTIAHYgcWsUWL8tCQ9lEq7u0RG4hH9rP5FyjYGTo/XIbn3b/133jk+pXaLh
tYIASiTd32CUmmjEU+wueBMp79cUFfCmgAV1jYfcATAR3YfW4DWkMaSlsE2yFrLe
VJzUOJjxRC/1gKWObmi+woHI1/R4DCV0G5LwIEn0ppUeezEcmQOGqzupsIrJYk+G
VlZiRlRwAxJXiGrA6iRmJ7AF4yKl//2RfCYIGERM/HHhPtdsK/98svtIhQayr5PJ
OuP4U0FZzUS2hQArbsXaw5Pi8f+Zs1jVijY0Vxi3oWeS1s9fGjDuduQZDnVh6sJm
nCAW8UT1A+9KAad1/ZwL6/mBVGJqiO0f/jXKX+JVj4sxP0EvdXFQlhgioGBasvTW
5UWSt6sdQuRvKZLFGXeQAsIWlbckgEWSVeyRMAbpn1hes/bLUkj5OoJ9lK7VcgWp
sapj9FMwV1MeHiN5W7UoDIu+Xn+d/MV1dUWePDCIUzOnlq2KlmJYzgITgbJimwPp
ZBa4x6cWs5ADTJI3JyCP/ftIp/qajgBklATl1OhMaFotBzhof6w5NhuceInEtOGg
lCYdzehdcXvUdGbiPfHpuhVLhkvyvqQ8Nnlkpe7S6MC5vqmjQHFC1tQtdiY5ygF2
ZdfVBj+k0BUEPPmEohmUAkzRkaWj7oTdveUJ0UKpTGN7oQ+JdGNZ8AdBUDpCwttN
CtKWRCaaTqfLSjiuRoJ8MMbY4WGAkye2U4n4Qal4ei3yCMPqeYVJPr9OitIQ18kv
mGZARP4FwQsBXnm3EzdcNT9TCSb8GZspVXo8b2xM5Gmgpm1PcGGtCe4P993wLNWl
RGzHId6cORH2vPVVf+bBREZhPu5IezEUxxoAmfpW14Pn4fgL6BmPGHiJ1+5LBzYt
sfYTXKDUjuqiWQXYWsEkvFIn855uFg6k6VVv+ofApN5VV3PT9z+HFHPLfqw7ReS9
RjTX1/057tQY3WXKXBRexLJyKSdh5vyT6c7fwtqVI9rhQ1bDxWos5VjFsVdV17pb
ZzSJJzzlOx3U8I5RUm5c0LP4LrsNo5jlCFFcCoaDf+lPm7B688LKyuWIhaIbMjMH
Ww+rl8HZGq0hM6J24TAfQLHIzWTcjuFTtoEoctO4i7YVpCt4kDLJ2vhsiaG7k5xi
GrZCyCYBs1d/eGB2TyaMD8uNb7yZWTpMGgY9rFJujWXvrpoFDJzgLrqNGcISAx8b
ikeMUBKFAauZNmCqTRfE7W+Lo1elOMhAN8g6B/+eYZD7B7KBpCEE+RrHwlzmvlGR
3uvuobgy27lg0hPcx1JDjkrPVoKVVjRdL7szdcdL+90qbgAwpQseLs54/KOp+Qoi
hjzp9Yu39xG/twhRk3bixqM/nDd5RppX6xkSL9gRsR4JPv+9QZbBpd2aKryv3FuA
rNoaFq7n+thXsSYrnGygv7o4B1hOwfimeJZ88eQnq8aAdVZlAJ68bWgtWOxLx59S
I4xKoy0S5e8ODWD901A6p8cd0Bca9JQxVeFqpHZPQCHD6qY5fdoIBbQe1k+WAy++
WFMHnKDYpZ9XGf0G54UtDVdKnXEKCN6719jW7yjlGhUqZ9C9PFIZDWFnGa9xMGOb
Y2k0e+w4w48HNn7MnaMv+pV80+AMBd0UzZ6Xc+rU9o2vgnINcebLJWnOBAyPIf4T
GwKmiPGMDK1Hs7aAn2+CqqH/b+PNOYOj64xMNV51yLKMViUOZkqNG50WbPDw6Vv2
r5jJfuD8gJUw6R8Lgcde3rYM5MN9iJ+hSm1hVq4ai8oNvmBKhPC9DZQDMtrFASxo
Jb95Zv4ezFvhWckSQjonCghImQrMzCFw2GeAbobnP+2Ij4vA+Kf6KTyfZ5AhU6ir
Q9ZhOxB1bWunYwrWLlbTEEYbIC/eGTy3TVVuLAIIsUopEXasl7pfJxi9RAED1Ulz
wPF51Rz8tFIBgq0sS5uDDz24TEAacDBxaze+yKZmyo1h26yxI7UqPOxJ+BmxZiUv
gJbgIvmHhcc43gz24KjiVE9ffdeoia/EZemeVq9ia/6yDL8HTpjxhKp63uWpGQfd
BeivwyzKrhKfCRdNSNEZZ4poAgpRCWlrO9NmcfPLTRLNVCYs4K7Q03NCF+jfM65B
28XpMSsSio/pTnRp09XMOw5mtz6OkCoAh1YzHPLsBKQHZmadHBpv89h5p+DMxgr4
bjaFhu1JfZuNR3JhMRzaV0lklkeVUhPHSkgWO2TwEPv6fql/v0wzCgqfRvd+LWcU
H6ntqhd4U/qBiG0ZhDhcrrPhirYs9yl8J4GVmsQInsa0K8hxfHnHVjTDrCJ7SHay
3pajfuN8ngrOOcCZMqBA30wIxYLrRpwdk/txoC47ocvXlkUM2RFS/cVBZhgCRqas
CHlrl7pEMVbDdrMu2qZYI76aiOCbed5j1PI0XZVFwG9IspqRO9kItDQPQ89Xe01H
vwJm6dZu43wpEa5xUdUk+us8wHowoNeBqfkIzoLMlDBwNBJflvSoE+NNic2yPhOV
LCCgh3P4v3xMPy5FluEw1X4QjKRBUnvqbErhwaRhALaqpZVCBCCPkwlicxyVEzmG
U6luFE55mF2dhesbv+37GMS4WdcxPvXnu74lDnj7i5AK0vt7dtm5TvvPwV1zUycV
zMIH8EiDbWBkK6BuLvcFlb2Ft01W1Sm7DyAfO5YeyoEyJc/TIBwyl1nREBoCbmYL
vwlFmiUmjuh3T3kTY3+4srRZHSDg3IHd5fqoc+J4y1zzRNA3RyIENnFYLwMC4bM6
/8Bt2+MXJJUa1dlHelNV5ZB9e9KH+d2gevx9YFL1R9RsU6s3GHouyba48oaHHDCd
LtAQSELo11Q4CaaeWyN+8CoAtHtFWqoj0bG1N1CNxV/l6hC58t7IFiy+YaEl9d+y
NWXKbskingJVAYJGnc69FVy35OkUMKpw284eS899TvBnhF8M5+mDD4mbhQgm1Pn6
Kqsep8xkWc40ex5ucvXaf41jDmsDUxqoIQ7W7ttGLOYIJ1H34Lq2/jREQy2egMV2
d1R/IRI5DRcS7+UKOtmmhmdeEHRwMjHipvKIuIFqy2yTybqqcYMJArVyj1stms1r
tPIIcjGcqzV8iY39Onl0dT/U5sPnFLyrREsqxo99JGYmVKi0NH9xvUJ7Ac4G35HB
XDFgxtIEXsiaB6KA52SDQzyr04ei2E6/XUKtk+aKY4ntAX5goteiBFeTMvZeXc9B
6wOSdMYn7NLTwrm38zxZHfRa4JU9vT4MWuAsMMLhSmRyZjKnZDZpEmKHCxEKqudN
UF7Shlk/eFS0V/ybhgfrTJH0bYl9zkNg+iBRO58/FsHDKRYNumESIPm/leEOm4eU
s74T1OkkC1T9KOxflMDnR+BjknVUSJ1ygOn5KQMKeWEqU6GyxPu+4F6sgaLhQtvW
s56BqEnFJ/45wCMio4RW8nk2MkNtJ/1ZVetcFDpChPdPNNGFMfZNMGxDDYDhU+RW
w7oyNLzGFBhsO1DRnG4Y4xYdFbvWJdaLFRD5LCBhsh8RdOzg7Q8/hXcqcAxpGlg3
eysW3Sqf0SawidN3dgzFlCO/EhK78sVAeBnKZxVrZXgDghgTf+hqpWXZt8LHL+EH
AYs8sTZ1NR1UNSxFY6OjFMS/hU9pm5bgnYPdqkluVjsMIYLRDhGfUPy94xTyTlXR
2ZqnffR7Us7mwCar5Dp4QdSnDAvXR8uqH3QvE37VRgm6/X0EY3fU1XBUS5tAMEI7
c2OyXSBeZbXJEdQL88vHVadvDuU3tHR45d/xHXskRD7IWX6FGOPPU7ulV5U9dDFs
QW3TuppQa5ng8ZwXzYyM51OhSdbl6j3YMTzGZAavFTKC1rqk9hS74liFK9tclFx1
8zZNB+2ficqo2Zp0Mkh4adz6C9O9CObU28dAaIbMy9bwbifP1Mc/ezL7mS/msdBC
bFppkH2qUATLfJKFVT0Ziexf6ipKs/lABvqBR/I0v/tqXMmbeBbRF/pxQ4vtqDUA
AS6Fjo6tzc9OnjpvjUrxU83FpQ8YycthklV8g2gi+rCn0nc/p8j1tta04AdYHcxP
p9uQ8OemJucndWvRua6psvDtMf35Eem6DSvNh24aWG97xjfCAGhaxWaGEZ1SHtVy
uJ4KExPKXvqxL1d2eGkv9FjHtg4RuYjZmKrJR0ztQG/zW6N+6sOG8JdiRaiR7ctG
YUqnX5frQtlLcKjvPZDHyiniJEJhKLsZipFt8azpcCl+kqNfYgjyfLiR0XS6HQbO
ExtjkQmdqYpeEzGeEJs05SGnQBHT8EnuTu3MPBgeUokaPoRlTO1NMmnfadDPnXTm
8ukj9Y0sVFsgt8VjGn7Xh9JvOL6Vf2zFYvxQVSRCFLduZaEUzC8BLotRGwVRr762
4ezxV3RqNoDgcNDpwARYLCgPzAZm+IrVYpAHqTkbbuZqm4uN185D1xNPmN8G9FtO
RP46qqFvaxfWvbJ1L31fitjr2ZjEjpyz5aO0siL0/m+UMy/oH7QJXbqQEDVq57HG
MbqcVhkjqgmWeLmUgIDXlKf5qG9d6r13Tx3tMR+vJrz1a0FWnPje3bWzPrTuGWr5
H537YL9TKsh1iZYWCl7F18A2SZcxt2olk1JnvGM6bqRlsW4dx+OdH7cimWoE/bPL
RPpso4gWcApmkiGyJw4WlpjhMWB4rlhcUBdnnK6W/W8kEAwrYQq7i15iiZ/4eqtW
Gha2/vTfI1FH+7fnEDaLJ+GHP91ua8y+pN8MYgonyJi6tPhuZw5StWXmriVivsWL
MrGssNQJK/LHJCZm4LS+w9DTcdqAQbgkK7gi053APfmht6MSFRO0zipHzzNr6RmO
iaIOS4rClkiZ8f9yGy7Z/T1vYVWdRyvq2FmPQwFSPhCP11C6lxvvtTxbPeivD9fK
EBbyGiVpk48LlPNQEIfqvKYc9s++0+FVaKgvPMiC1atXI+3q6eagmJpEzXJT1ZLj
z0vvEV1oNaz/nr0tiztxtjXDL5rBErFQQQpRN7IgE7yeC3KyyxGJ0mi4PTPpswPB
F3g7mRGkTReH3cvTi6aTCDAblAKHT9BKM4PhE4D845MT8wBftLBiFhojnnujNmiw
AL50gvkmOl1Lq3H1iuaOGYUK8uusioU7w+YIsTrjqS9tnent9+AybLcRggiyktWb
I92CB0NPwXh7XEURvkCUoc0OjgHgSlmcOaD7DEHnu9g/62FUBLh3jV3cxY0ZT23u
EYlieULpBfNR5PuT0A2QERDjKtPONEMTAGMk/KhH2cECPNoMWLbzWGhJLHEESuWY
o3QrJwMf2eGG1nA1BtawM3LZRMUtC1aqjoQWT0ezmHuwQUywyswhf+QvjBkCr4x8
4Zx9mDCz9TQkQdZRQ2pgJ71gD3HlpnZwYBbsJzORxzjxQq+nkffd1oeiIgpgLcrL
Txm3OI/Ko6w4gkdIkvpvGSrmqdfucIh3lp1UguBsKiFktyNoSIuNowGz51i39JGM
u/mwMl5B/TmJLWVpmBL6Kh3gaCHdN1zLfwiSF5qA9Rm5atXZj2YDNZzehjAImhnr
IJcEkcRPuogaP328jBbTc5JAJTIh6WH8FMcrfBlEymlh4NHilpc4nEb0AEecGD8m
55DpNwqseboIG5/6hcxLc8S5NpqhwIpaWh5U6o9NH/1c9HVS/8rVd45ghfobZ6k/
XIhhn2zTGbdZhhBfvq0hSL791fEkLhFBmIpJizqxMCHQ22uPgq1HkIEsfDyJeaFt
zOoYjoloYuSJLAZ8TUF9ahbWpgrhUsl4Ho1Z2Ikj36ShjhamaSrcbk+HshtaUlyL
CAYERSpP1mvgQK+ngp0WGluEExVLOiz67eD88I4Kg2lDVscu9lunGDyL2i9Us6Mh
h8O6Y/E6gEVS0Lq0WsbTg5HRcl8v7nAezQQHWXh+u4q/6R8RHLxmiYVK6drUR2Or
mfybBccni44hNpwZSPHzlzTPLcExRngsxRs02zyNAhc6unc28DqNXT41kGCM7jl+
OcH5VDaUSD0WVcUogsqgNQ==
`pragma protect end_protected
