��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�GN�Џ	�UQ@�m좙�m�/�"�^\��>�k��lf}�˄�	���b�g�Ծ6CζZ0��J#T����=���gn��~�_0&l	���/��D$�ܔ��������C�̡k_�����!S[�f������Ϳi��Q��t�d�P�2BE�%kD�T+�u61���9�h��g����4��Ex�M�SO�K�N�Y�$�y��N�f0VWJ[Sl{�:�2	��{;�;�<�7y��ŗ��)h�iZ��@����)*�em��I��ɩz@y�\.����E���� �*�� �5�VRT�-����F�0
Dn�	� F҅�'^�_����H�:��j�Lh/�B���Gd���r���d�\���0���@x�˰3����bpb�)
�ȡ��<��d���
����_�S�@��?�%�E��u����26�D��1~�yc�OI��E"��F �ju��v�������$���J��/_��XtA��_8����`v�1���q4[AIʛ)���0f�	Z*��D1���J�>�F%�0�� "�U����Z=i���E���>����.�;�4�a���(P���n��@'���i +&�3�Ţ��_��@�rxSSp�� w��҄�vߥvT\p����;ܕ\���:���FU�O�a��4��&�a�?�\$�$�n�8��t�:%`��K+�����1����yoR�p�X�<K-��g� ����`r��>/P�$E��Sh� �����ӱ�ur/HI�df���f)�.؟Gt�W��޸i����u�W���N���1M�m�R;+���7
R�^Jf��i	_�M��L��	�}GM;�"���H�����!���?ѡ4����Ʌ�B�n��Ϟ@��H�H��xXq�շ��#t$9�-���>+���%`��&s}f���
���C `U�������;[#��w^����u��.��P�o�a	�H��gt�Q�E�JJ>���h	1 �2)�7F��Y?�xȢbӈܲ2J��Mw1�z�������v�|���[�6����Ϻ���3Y.Vxd�wu��٬�@C�%�p'��=LL�IU�����m��G���L~D2�zvd=�_Il1eH��<�
�����ܯ��OF���K��+P�9O	$+;'��#��[�]9��7K>Hi�� !}%��t��RuF��Ѷm��N���l)X$��\���Y�=��K��g��OHV=��xܨ+���tm��fK��k���p�1
���h��8�����<�2� ~}���CY9x]R����?|�d�ќ%�yܛ�hw��&)B�,M�<O�/��F�����Q: u8���ٹ㰎����$W�3���o�HQ+X�p��/+ֈ$�g��}Ņ�]�����)�g�qZi��ڲG]^/��N�t����w⼍_H��ýV?_�D��|�ʳ.u��M@+���?Q�e~h.�i4&�X��%�����*Ėn��slR	����I���ϼIk��#��-���N��"��0*�'���4L����ھ�\넼�tdv�#X����$e���7�|���:�d˃�˂[���9��R������}�q��ͯR�����|���~�c�7nT\^F� M���^�e��DF{Sj�A�B�1pLؐ�Ӝ$$<~���e?]V'�pe2o��|%��l�iC����$r���*��M��=��;�����fQ���9�ٕ�4?�hה�����gY���^>�����1KQ0/�J����Ŕ�*�U"�m��<Go\�C���!�pp���N��a*���f�sai
����VqNhU���}ҋ,
'�?��q�D�g�<���XUٓ���|K?[CK�=o��B���~�M�
SU\�0�k9_Su�z^��ؤmbl�rk��*Rl�Є��[���x��_�s c��؆-/�~{������2�]���|��C��.���R�d��_@UB�����=(�䶷b��Z1��X���Ӳgҍ0nBs���Dgf]���=ߋ����=�i�Z:���QZx�Qd��ջq��o�=6�ʻ��,5ZBw���iu��{i�е.�o3cucR���-���KL=�|�G���@p)��?�8�u;�f���S��U��n����xH�i|'�C�Bz�ab*@O����d�V?�E�H��3�6PYL:}�Q��)�2�
�n�N�I�%�uyR�CpT�r(�}�3��%�����.euW"d���5���*���8I��6�k��Vsߓ�?��S��b2��>�<=pZhq묤f�Z���}���=!}>��S�״Ȉ{7����|�f	\�Md�SO��TxjR��b�	YK�(�׏O�"���$�������}�)7���뀛��ڕ�5�,��ZV�Q#��|�)�1��7�-��D'����9 +�K�����|�ɘW��Ԍ%�
�j��A���uUJy�8[�-�z�-G�u�S��0�1�F� kIZ���ZZ���|{�]�6��-s ���c��o];�����k��2u� }f_���|t�h>[!&!�"��H�C�e��ͤ�|�9c�F�B\��]y��r�.�!�DӇ�^hl�ÍZ�#n;��=�?���Ve	p4�?�R�qT�B��V�-��'����낟#���] ��Adp"A������*i�:JT�,�xq�٢�&<�X|�,�G�g~*�]J�R��:F�l��Y����=��i,�*�z-�� �2=M+Y0��,j1��KTC�O��IZ@M�:���������7IP�r�}���Hw�MZ�Z:�5j�M�:�B~4:(M�;�^
����W�j���CI�n O����f�7��×v�@53�j�dA����~�E��0��K�?-c�.?
8�n��P��=-��"+��c�Ae��'������΅y>��+�/i$��ʚ�#.��`�;7����%�@#�Af�ݫWZ�nq��t}W>b�)��ބJ_�b�͑CL��Xy��YykOK|am񠪒PM�[LpF9�b��@�j�-Or����׍Q��pZl�T
�?�X|ڈ(Av���ğ�B�0lG��6!����S>�D��I����-Q#[Q3�%�M��~���2/���3��b�1�08���z���Őj��6��Z܂�l$o�� =���_92A<�n2b�>���FU�Q'��V�%�$}�^��[��Ǽ?�QW���Ĥ��yE��tXV`cRG�ߚ�J+���nȌ�(�x�@@�E�T�����v{���d?XPLб�!(3Z����>,7�߈ ��%r�ԿCﬓG���4�����ñ��a�t�F����=���Nј���bA��0^m��bm.!O�����T�W�����	3�*<9�/h�����و�o��P�(W��隀>�.�� �e��څ@���V�G����'��S�?�*O���X$�D�%6�P���"ˆ"����V8�_����u��51
wF�?sZ7�%/rԗ+���#�B��&�RI��$�
 ؚ����a]�Vuz���%�_���	�1��3��d��ǰ)N��&�-ƨv�`�Y%7�$5SR�?��6�h=^���o-I�=�c*0��f".t�sZC��!������eQg�|�t���M�x7,t?%�S]�R�>|�Ń��66^�������n���:,�\�K�hsZa ��N��e%@n�b�5���w�,Jb��C�9_�f�͒��֌�Xg����ט�ss��"6���L��C��B}2,n�F6ׇ>9��Ȥȍ�ԯw�IIov��^�dR���2�z`ꂨW�Υ#kA��t�0A��ى�����x}�f.؛����E	�SOZ�+E���8`�9=~������}������+��8l0��.b��l�ر�$F�������<z�K�ߙ���&ʆ��%R�Gzwj0D�G�C�����
�t�x�ʖ%Z�� #��R̷��b�4���bnpZ�j<{�ckz�dPuDGk;��éq�������*���D0�z&���=�ե0�W�L���kh����\�E��n��C�g����\�r�(���:a
�p��/.4w�k_vM�H�C��i��y!Z�F���n�Vgw�*�i�K�z�{�����.�'2/�#�ʃ6��ܚ�ͪ�o"J\�a�T���n�t$����)���n���������=|;Za�T�29���&C�z%��*�"���� es���5��Q�DiX=�\�nqLh��h�.H6(m;@���Jm��k	7�!b��W�noj8L^�z��ܬ1�/�C���W�(��]��h�K��Y]������!���&�`8�`��Wb����Z����KÎ;��]��B<]�:~ir�*+��=���G΂�5V�h��(�`+�e���ʀ*"R {�WG����� ��ܑuAV��-�n8����
u0^h�gMJ��;|�)�fA�=Hl�J�i����?�ò���Deu#��#l�ED��r����i~iS<��^��ƞ��ڕ���8�d
�E?�ġ��
�v�8TA^�j�x����?r�A3�tקi�1���!��8 ��<�>=I��Ͱ���Q��۴,��_i)p�8d����-"�̌*��8-?"�AC�@U�h�[Z�/ȥ�2��`��è�����D��p�;1���м�<�'����7��ƿ��|�.Y�q
5���S�[�L�Z"��ɟ\��g�tS�*��vy�'K��l;��׋p��?��osFYQ�r^���
'2v:��#L�%�wAk
��~RN
J�6��$(W_�I/.Ա#�c��L<Ve����&�L6���&	����X��I��9H�ZU/>_B;,w̞
o��ը���vo�� 0My�'-�zt�I7�&A:r��������֚�� �Yo�fc7*𛳉ۏZ�߲M�@��8�Pb` V ����T�z�[����~J4b{,��X'C��幖��3����W����'�tPc�;������u,��Z���m�w*�1��E_��4���,0SI1W-H6��ǡF�Gt]jX�"3na;;EGPr�8IO/4��Zn�����A�\��$'j��ɞ�/��}9_d!����	|B���&��'��ؘ;t��z_�۹b�~�o�dʠ9�F
��N��òZ0@��v�g)��J�Yp��O�\0�	t�����$��*^W��a"/cM�w������_aL/�,|qbw�����%?���3a}�"4�"yk�e���5hQ� P�W����}�1��=IΚ�U� �f&D�sE2�쌾��,~���7��t��a��Y���}�f@�7!_?���+\00��P�Zd?@��H�)���ՈQK�C��c�5Zݢ�C�_>��E �o���m통��<Br�����ד����T���LQ�G4����<#{�7{#���3߂�~��p8�����+�r �Y) ˨������\"U*h��S'�{�:������<��j�'E�Ι�z,_@��c�w����6�ǩ;�M�(����W���ʒFٹ�EtI�Mj�l}��hݦR���Fd@�������Sz���q���������t��>��c��(�;���~���&2F��4,Z��q����r���~�>�4$Ay� ��	x��z�Xl2��t�L��O	/K����B֨�X^�v�G�%Jy �OT�py0˪#��'�Y�%b�~�($3\�R;�3d[h�lh*��y��/�jo���K8 �Ƅ]u�!�@��l�P �?��_�M��evD��$m��L���_�������wU�!G��1ԕW��$����GP)�`0B��*�%`���¼փ9�3&^�/�ZA�G�ٍ�2p�6�'�p .�;��
)��|�(�pl&�����:��:�%�:ڔC2���Uo,B�\KJ��eT�����]�cUfK��<��dV<��� ��M�h��,[$�����9��x>�V]9H3�3�ꇼ*���,�����ke�����XCKv��W��i���a�0up&���W94(s�����J+V�x�{���X|�6��r�3�m�]-��=��|l�Nh*��9d�Ĉ����6#�����Z#����b�<x�=ـ���7"��]+�2�`� �fe�2̜�ߺ�+f�^�.){�AZ�̜���_� JE�th]��`�i�q�����=�B��c��뜆�ϵ�J�l�����*^�_qK��Cˉ*L�R˱v���&��H[��X��qv,�Z�WYa���k�S�Q�h�n�-�UP��Kk[����S��G92��o�D��P9��bEM��\��E�:�L�;u��8j
�Hqn�F;�ډ4'.|6�P�BFk��r�D�����)��ɨ ����~B�.��1k(>)��1��F�`���ƛLY_>�UN����	%�$]o�����4��x���L�� M�Y�s��F\C��ۓ�����յ��Y���Ϫb���Q{�j�9epF��h�"��?k~��w�O;av��ۏ�^�V�Lv�*����DϣT�B�n}��]��j십�k�n6��*�1��
s`�{����X>���L�����%���6��^�!��=v���w���������y��uZ�ꖵa�q�/ �R�
y=i=��d����e4;�`��ίVD+����1QRє�S�5FU[F�x�����r�Vd	z�|x:J
T�K��m�V-E|��+-��T@PB�כ�>?uI��z��F1O�?�-a?��Tu�A�*�2n�$�Pȏ;���7i�7t��~�}}��mF$ȳ�f�(��Ay�r���;8�r"�� �
%>���-�$���$�{�{Ɨ��G޺k;Q	%/���z˵F$�,�`3���
+�Ǒ���� f��p�0��6<�9����aj�ɌI?&���f쐦e�ԃ���J��V�KAA���
'��k��T�&z���+C�a�^Ϛ!h�'���nZ���RՂ�t�:+<,�_1�
�/��υ�>)&�%��n&I5{M�
����V���	��q��&6A��kMKY" `yƭ����ֱƎ�W\J3��S�B�����_�����VS�	�=�Pfu������r*�8F?��e:��.��cW妌#~n�q�:��D�̪+#�P�~�3�ڏE@Rb�G��p[�8��>:5�p]2{�o$;ⷛ�~�C�r7������o4�P�Jm !<=�@b��]���Q���Z�=��i� �@��Y]���[n�`r�0dU�bu�
��D�W��J5|��{�.�ݩ�K[��_�BU�^38���B�1���MgN��2�V^k�ի*�Q]~����-��֒�X8�@�q��:�2�'�
9āoc�R�z���!�
l��ee�s�;�}+�KhP%��̰~�޲co�����Q~�]S��}2�sq�Lm��78n��l�D�Q��Y��,w �1�0b��Ll#��ȧ�͚�����i��)S�DA*���gStW�9���YBBI�Ihw{>P_�r�z��B�_�W:X]7`K�m��V4֋e�u���FP��n�?sk��v�HM�X�`���p��,��U!�� �g-Q{f��Ϻ?dS+^���*��u.������4=u
4�s�8�4}C��v܍�a>���������/�у�ȸ%�ƛn�LCU��DXxjLC��Wa(5�R�q���c����+T(�ntE�a�@A�������h����$ IX��@k�+`�� ڪ���!��9��G������r���^��-�!�N�1����O�葈J�K��.�//��(�7\�9[\e���H$��� �-�)�wo��[��(��%�X]㚓���qĐQ�D�0������F�t�>v�:�K�_�9�M�:��(��P\�5+�4?5OU�o�t+b����T�=S}�>Ub�e�,��3�ы�2���.�J[$ 4T�& �Fm��bv�Hm����	/+0)>����L�R�P��h���<O�l��T�"d���YQ{eh��\a��ɠ׹�
d"
>l�h��u�m\/N��a�d� ٚ�-g��È۵{sA��+R �D����o�E��l N@�z���N&��	������`UxT�5���{ϻ�7s'+�y�A�s@0�f�d_@�=ܠ�Hl�GX�,EPԾH�����x
�ג1�8CInAZ�ko��g��NqI���Z̰���{|�|�Ƃ)��`"��pw�^/�s��Nƍĸ�3��[E��.��2Ү�۝�i�h��3�,�	Z��'�.cu�Rˍ;�:\�!Ji��
�s�i2�i��{Ͻ�N'1!m����U�^u��X��6mj����?�G�	���vz�܈�[浈l
(t?�zgm�3L���RS�n����H>���p�����D#�/�����+�S�[](<ªm׮~��z������*ry��+"߫�)���W����x����$b�@s?�Oa7н�"gvS;���]ӟ��ف|��*�Tǅz�v��C.�����W��X����� ?��Zf2{�AӴ����:�(�Ih��E�MJ��jV[Q�1�je����p/���,�?C����Y�u��C�tT%"n]N(�q~�iٿ�����:��{�@�I�>La>jК���#�$���,xFq����,�w����*.�/���o�4���$n��NnM��0�(OLK���Qj����8r��:]���HC	�������< ����W�O�b_됆��Drd�}�9���!�{�������o�.9#�ÏU��r<>��y���.���k�/=��pd��D6t�q^���g'�>7:����eQ�f�j�ӬyT�(����3�Jk����e,��љxw@o�Ph#�&|����i��Р�c �w�D��0G1��ʲw��E����Wё$$�h���q`sP?�(�NUz��lg�tD�b��eJ��l���]�&�?�^ q~�sQ�^�S��E�֢q���W*�V�V�j՞��!��,8���6�H(�"��0h� �38�<�v*NX�UU��D���i��	 ?3��';�9���u�ֶ͢`�g�W���ծ u۹��_v�u1��P����4V8���P��s�Iʜ[��N����g宛��%�=;{ya�O$���1F�4��N\h�֩���.����}(�F��(��H��yk�#��~���陧2ʍ���h���s5 U$���b䂸x��i�"Lo��ǘȾE�Ŧy�n�`* �C,��0����	���rf�K�b��<�v��,��R�⨫p�Dc������'fDw�|M�)�l����׫��pV��D�]}����|����@ne�}y� �^>�.�߸�p�Z�CC}'-)�5��+�b{2����/����I�����)[DA
g�S��zW�eyk�2Q�������W��&���Q�]w�?����	ڲ�j�n�G4�6z���N)V�����Ty_�t����dpQB�-񞧭����Jր��_/E���_A՗�����̛e2����iX0�Q�sj&����<x�S�lY�S��6�p���9.� )@i��KtF?�m�Cn��Ҫ��*Jrj�����y)�H��f)O���ܪ�O$G�MJ���"��j!��׃��d�[�fBp�2� _<��e����7�)K�kЬ�}�󬫻��k��F�o�2�)i�ʷ���k=��+�s<?�_�������O��py�R{F��X�QWrG�����^����C�Ȼ����"C�c���V� ��N<�.Z%���B�^?��m��dTj&GG7	��|�l�^
�R����ڃ��u~��R�\?�T��[�j$�1 .4�1E]�p*��i����2켁�� ��$���D8��b�
�������%����S��v����F��g�f�.]�]�.������
�畅�f�lg!,MLRn��
2TI�?��+ϫ%���L��h㮂�
����ౢ���#�^H��
H�S�;�nklW鴴_���4�+��
ʒ�m����^~�q��j�a���˧��\��*)��f�@▁�_�^�����n���B���0�:.>ؕ��JP�&�GS<uPN�$>��F�f�l�m���8Ӹ�)�s?�T[.��&�8CN�n.Z[�f͝��9t�.�q��|�j>ۛ��=J��rb\�<��F��ݺo�]!^!^U-�eu�@x+
Sݠo/)z�����|f?����)]���V^�D�P�ǄzZ!�;��HUCB�4�a>'�r�g���K�^Ou!�Sx�$gEWC=,�	�vm�1[C6.f:M!-W����0� M��倪Q���,!��A�#��s���c:~�:����e�ʫ����&��ao7]^�O�n���z�����NQ���4�ȑ-FW`]xL���M��G3����g|���Gۡa/�X-�_�b	Y?>NEA�-~����wx9��s[��R_�L�p5.��N�s�(����[=�e&}y��|W�0���'���Cs/�q�Z*�*&��].��W T�� ���j�Cү~�?���P?~�V�EUV'>�3F�1lhT˂��c�2ә�?~��̘F�3J���)�QA:l�L�NcO�a�-N�a�_̵� 64.i��Ծ�����ǆ�c��>S� ޳��s��㮼7�1��9JC,�#]J(F�� :��{����BB_|�k�O r�q q,0�VKw���(h��bs���C�E(�߻�;���r��D��p�'���<]���җ I�-LH�g�=���p w�"6�s�2�����2 ^ F�˧�B���A��ٗ5/�$�v�r���+11���<M�KD��ԭ%u�`���{���I�s����c:2	�F ]T
��a�����Li��gj���K�w����9�v���������j�9U��#Jd�Un���}����6�!��\:����W�⃖��k���')�~,�$u���F��r�k�^��M:��OI�g/b]҃%��.�w�#�lTtE�,�,<]��/au����xn9k���HY�9ٕ��ΐ�34\�����_}�v^��[����(��9�`>�	�#m��� �̇�vb�h��E�r��+G���x��^�/�XЙ.��,]��b��ʾ��)�h<H5��Ɓ�V�C��]\���xO�9p��d�����,��i?iw�0�ݷ �U����ǬX����쟽q�&�Y��-0��{#\�<g�8IӰJ, \�n�H���uXr�y'%c��Ư�1��e��.t�ls^^����r�J�����-��:2�=jDGf�M4�g
�ݚ�%, �iT@���֕c�#>i�uE2��؃��4����,�ĭ�Q�Nabԙ�����-�%�v�1��V��^w��B	��n�d��F ��J`�RUՐ��F�t�9�U��b��,�N�-xe�����j;)��h������b�\w:�B���� ƌVI���[C������ZЬą=���J�i�z8�?�[�#|�8r�Ez��ɟ�t"�%b#�0=d�gql�H�`���ڼ���,	P�M��ǋ*���xj�N/��=Z�h�'�n&h[�~��WY̆�#�?@'�j�*�#g2�.p��������7��f�w3���y����r��ڏ\�5<��imA>xt�`$7�M�hy��d��P�_�L��~c[��#a�[��jo*u���ݵ��K5G-�R(��b��{����)�ɓR�]l���3�_���JFW0���q��	��!�m3�+�9'2��E��0��!+�$��h���̝�r�2��Չ�����H��"e���,�"Z
(~����+�c��G�?�W-k�*h�F6n��� VUZ%��ꞣS�ɠ�y�:�� ��'�.��u@�G
�H�N�ڭj|���D5��l�9ȜM"m�~]��]\݇��k�J�vA&�Տ̗*����	.:��;���@5�JF#��UzT��-�\t���_WM�[&S��E!w9<�)n'�阄����%����p���q�!���$שּׁi��)�j��@ve@�>x�� ��9#p�F�3r_���JF|��%��Ǆ*����l,��!����S�LC~��)�����2ͦ�o<�0�m	:�i��ȨrH�_m���.y��P/��\����4����5n-�»����; �U�*�A�����y�����^�~�u�`M��e��掤w&��~ʕB��(G�~� >�D�1� S�}�եt��|�ƾ� /`9�t��Ţ��0�����/k�3t�`��i�� ��T���s6� ��L-];�R^�%�_%�!>!��~�J۲f\�f1�s�GT>T�%gʘU+(�q��'S@t��ή]��TE��c߿��>%��a����A_;