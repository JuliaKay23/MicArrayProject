-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rX7uTd4mNHPcHwkp+aqLL4swaQbVWDhdQpnqv+Xb2+wrVavwOos6UsZh/XzVCnBaCyKkukyOUnFv
lHHjKBx73gsef8b7FWz5sIqwfOyteSh2IyeY7Cv0DSZl29zVRPAxu59o3DzsFUbRsvGwTCdfytkJ
rsfYke9MqRpxddcHJRXC9yGV6VDj6u/BEOjcUg3wU2cRp7fzgOsS1+FtxXqDQHPWiYKwQ63+5EiC
BPi09P3806QdF1fS+wVKvb0eK88TzKJ9j5+Etf7oy1TwfcFGn+nFuWOu2o8Eq1GsO4U+0xRD7TwB
18xuRYMKfYlCPF8K+tzuMtRoyKJPklLWR7bB4w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7296)
`protect data_block
SBa+/m/XYaKbIcA091kzwK3l5geQBvKndaLQBf5z3LbjslVX8Hkzhk9BoRQRiMUuuoHYnseCG3Vo
MH2rU3hdUQuk+MrduWhQSOa5fp97rNZ070VD1VivpGdOV6DiVKl1jC3LvC0sdw9GUowMs0TBS5D2
qnN6TAyk5OtFFRdwTF5dDLmcttOK/zpaEEoYn6LzokKPie75BrVckpbC8z6eW8tQaBDb2SfogAV8
wh4przMmoGDt50/QpXb+7rGiDG5QlHJHoExxF4zeypuvYpSghq1GeKjHpECMwCl2hW4KKTiIJ/Fs
DYIKepjkR+7CWl6MUzdxEkU7pdUgNs5O6dxIs0U5j3eWsgn10e7F/VkCWoeOd4YEevosMl1dzNm+
q0wleObj83qXsdK25yiuWPbc6hh8HkBZjMRdyDifUEMZBLyFcLPUvX9IDZNzxRDg0m6q9GV4ZaQl
JxgbIaYvCRvA/fjBDuW5revtC+1K2RJ3qqAhNnXuksRcS8zrKg5lTRlFvnQCN6EFvpiQSgvVCHAV
bCjrvWIbW8R1Pau7bamSBri5liJNXYLvU/VQ94uyeLD8iYn1FM2Bm0tFUSfF84B++S5Qqjdsny+b
WjL/OxUwbnbHoBcAlTJCFPAKFlQhQpGb6bBtxMq9sXMrD4z8MxhtNX2VwhtGUVbZkUyIesTmGPKO
5MXmtKpjr6BxiWhcq+/JxYH/Ozm2vYEhIkJCA4I/AchGpQ0IEiOWBE6QYA9Y/+I+d01S3lCAzQQN
VeKJ6P65aWSACXsHxRC5grKn991fPNSd8POOMD/BMqbA9nHBAcK0HCMrT5R+cwfdPhh1LRALOwT/
kmwx0hwahEazNqGm+IRoUXGGLZikEJrgYW+CqZpV+SpQmbOJ4zsGjUXoDXnVMzN+eDtgxjduTIa1
A37ITIXVRD4kALFs5aWTuf+T/STCwVVGOu6v2YfkquGOF1/A1DpsC4iSw52b12h689dcfChMyBHT
mMbW5mGIH6C6WFBbM52Xh0hz2lKwceO59uNpcUr3WrwTuvxLOllkUuLB7rCTPvRGcUjCQeTFhIVv
sL37YfCDPO3MfAaEQwcSjNxveBGvwGO8bzlATrHygbkQeXgsN3Xj+DeRBFV85DyB/Yx+wQJ56Hes
TtTBeFn313f1jhw77+fNVAlZXrAiE05CxJuQ8+gVEYKsPyaY6z56mLgSi6irVMo7ds7eip5d+bhR
gQx4cr/p2Xq19YMEg6SeTpLDY5fGDRO0VuSMPnRlBhf2q1llAxChvjqVSH5NqwSoCaxayy9sVqqp
WxmMhJXOMSRpJWZsE31cRgEMlgRxkTRKtsoMMxB0xNf4iPYsI4ZPthSYoUQq+LAo1a0aEgUYn3ku
N2olcOBderm9gI3xgnRo2V9glSgRlTDMfDJmSSaMcPeJ3vIcIHHuHxd8cYMaKA7T8vxKQoAz4qI9
++TGxMeqPcrPM9Km4+W7ttzE8mc/vzRrsJlMhiHGpdsSss6UtUtk5YK4Y1W0oFxzDBPCuV8W4oNS
TmJAT60wrzug6zjFRVh7PqtF5UfgHpnXH08fjWyqdG/tce4fhTy9GhGWJ5SkVTie+FWp7o9eTZlo
UwKBUJA5VYKt+rKy1LVV9OSKb7ikDC2AUFt/MUfBXdp5ancX0OS9sHivCSfXeBWyEWFeG5N2tjI7
PfvyGcfAkLMLGs6N3G6XRfLbb+MXDEjvnWiRun9MPdJ+lZY/CrLeEiXrrvBjZdghjMCgUIy3ArtK
oQcQh6TrLtfOS7Alj8NKHkBF+1WW5zX4OAvejWyDFpSy/p99cjsNeJW3K6N3fx2gFV+f++F0/jjI
3TIY8eIBiF2Bz7oTEFJYsIGwEm2T37mcc8uF34NE37Kl/1LE0VmtwZgcOPOSGH96+HAq8yNb0RBo
2/4+jBTZPmDW4M6SjQMieAhhxEwgE0MCrCm6avQSvSRtcJwATRsrvuKwJtPIUCCAK+gCgjHCGNYS
WW7zh6SwRTEQBh8kZO6+YFdg4dWyXMYRio+0+DsSF7/f6N3BjVNZfBaLkCkc3/hZz7IOgaZFwOYH
2XV4woFXUbdOHZLH+DVcufFKekQB50kaS12moB/eHlKLdQK9QbrruZfEEbM8FhvLOunUYq5RfjmL
AF8d8FlCDnd+kXh3hLi4AgPBcUTj0hiBZbvhgeDtFCm/QfJhw24t+SZQdRLZrak7VgiRouoXICiK
UarFrH/d6kIVxzj3qDfOeOqe58tNSD9E+OVX+/oPw+jXCyNu6H9earJpZYf01BHnz3bXfpogsZQQ
w5cjZ48LHnf5P5RTdyz4okDiNVw+JPEePcpA+PNjhnOsKhYTu3JhfhSqaD3FSOIf+9US9HCPbCH5
gazNOOTj1A9eneS9xVze3erl6R49Mx4vyhYnujTTTRPH2Ib/8df7jnLf42qIZ3oM9uyzk3hEguwA
HvnqY51lhslN+kiZk0uOMbMHb4V0FjR619dVxDCZHZZtP+dajfbJQn5oVLDXFv9kiRv70euIaaAF
u8/7EejvIA4s2EIpbXT5y5zmhcK2BLzlSGbLu2Yi51HgG6SGu/ZjGBCzib46czCnQ04WKJCR3TrB
2KrBzUNWkOw+eozLjWIti4arKIbtQXPE31QGaVLenAFk4XNS4xWBAhKl3JsfwgfRTsRPs03/JVQl
rdm6/RdYn6bV/2aoAIlIwmU9zyCgtCeHz/I988+6XWMfRwyfla18Efy679cGRycUOCzVjBCNGUwf
itEnNqXmdmoI/auJSVyEKfBMHgHjc9X5aX1BWxtSxg8nAZwcVurp647CtLfLrTLm2MhUvoRNPq+8
MlWiqBd9ySwW9uuNWXILWTO24iEZYucNHPfwG2WMCvUE0C7qUUUjLNPgHosB8Snb6gdXFKKtaKlJ
5FF3QHvv6qJOS2rN0GOGC8T6plTc5ouuJhLvCmZA99kvqv/RMM1X0rHRjtLDFrtMviC+gmngIFvE
P4lD/InlzXUlpTGTv0Vq3JUM3g9sLlCCBJnRdzR8nneXageztyfkFc9YcIAkmCCnKl5RgVSTaNMy
0oIGH380NT+uyTpFHvXjW2F07+OiVX/ui0Pb/PZX4Fi8i0ea12u2Goq06kBUcJ708vv5pfzYTXcF
xnncbdCF3siuA86h32+ZtMoeU33j0GoLHuVrpKcmzd6N8yCuG/jswPQYuDryPfSYDg32wQWiMtDG
wciDIwuZ7TDcPiU3FAHwannwVoIW+uDmi6l9vcp9556t/3ux3nXDiCUNOMCNA+TXf1hK7zKWa96x
Id9rrPUPmlVZnqwZHfQAnDR2JFB5zvb+do35ULQNbeOJZ/9M3+YDDdnR/vMYmRVnecIYGKuaafg/
f9r9UXE7xafT7QACqB5x+dM83CiiKhwTfj+SHrWSU+WohGjzBc9Kp/+l1+7WxNOMiOCr2BfDYBSM
yEusuFrOWSOAIWEkUdWtO0CsdgDMgFHzQd/AtDzowRcB9DzcRveYTfd233qYCiwYyav+gkl1N03s
VS9k77QkxtHxvSvuL2ZucjDCMV3ACi9Lvrxb8k+qZSwIDTv2jUe3xM6RLVOXrmjU423MY0QHvpLK
iZipba3m8CVYweIOe1OlsUc7iiCu7ZaO525mBp0lXEM37hHA9pXWwYaGigOx8rUCafeFdNQWxTWJ
1kRZz5Pyw9jPvVKASocs5lU6KnI0pTcnMIjSkKNkaIRNl0lhy0YfdP6XHZX74sQTRtUhHhgD03++
7lTi41kcN2rt1QFyRnfRpPhPytxE2sBDCctL1cFwqy2qqfT0sSkKYf9t39AqxthGn6g1P+bHZotJ
09GugyIl+TKwrjg2114XkoF4lnsINFH1acWs0Kee7HUDaeqdb4IpykYlX3QT/P2nFTOYsUp4Kuhe
eCklI9i3af00Hc4/siENYibPcvLWpIvb3SkagyxdDZxk7fY1Q8hpQZC2KEzymCBdc4/E2BnKWOXr
1p1JdVnCGk1Y4ra9IBN+R1V6p8GDUu0tKFexn+cFU+SLjIv+vYyHlyEks3W1xg5/Dhu4OtABBrAc
M1RsH6LmtBt9+1/zU4EGGbr61RccMkrJtZ7w0QVkSLp655Z33YFCkYETHz/t1t6YFtsrDG4AVmWM
2xMUNvDiLq65t2QTDVfZ9wPNVibbnrJRN+gslQF6HvNsCIedUQngZEtWwhw8w8aBpTaBIg/2ojAm
ygMRFRyZjd0piNSQKaUV5hn8e1qQhLPNM2U+tGVSJSO0f/HNRneM1c5srN2cWKsuTctn0GZgt1Vf
33nCSWIqdeJNpdsrtm13l+4KnxEWUpSbZDqoRI9BoCIFCxm/hv4138/HKqy40qtlH073UbKOXo84
BKVV4IU3yfTNJ5k1NfuR60N6BDayhBnUinAG9jV0aE77JYvOR8Nh85TXvi8PT4Pac5cnhYwqI34m
nYhIL4F4qs+EYtrlCjf1H4h0LniLrBkYSx2ruJm8A+I8aX4WswdckqlwKFB2+Pavrk59QT6Pw4og
5rsfSlZf402wUO1WJGKfAmqcAlWCksOH7uap3BryBbkhMhayVVYLnGcXbuV/w+8Nd0zOt0Osn8Jp
eHXyfSdG/9vZqyasyc4yCv8ZI/7KwD2+N85U79QWcMKucchol/gZDjNuxqLKYR7TLPh3Ys2BN/fG
Qwzy4J9bHSJ/Yl69w5gw+b9Gepq3xeFLodN1nz6QjLxvxo0GMXLioAuuxYvp1KQqA/Qq9LvbvRoq
UCGHt8/sZZvQfFNA8i8747MjVh8EwtoZsaNOSfL580gECZJ6gb0UptP0xyQB/ctAFVQjhZCNICS2
sczfND7BSpXyhnOfRky5SRHwmSDSTffUxLOGUVfAXbFCaH2qP8WXcWgN/S9t4k6IA1gefZke5r1z
ZtIrPzPHSvKB1yFym2rqRuXCn114JbOK3sPn9k83YT2+r+rzGXB27ttcG+bnuSB7S7CusR2pIyEi
jPIyspxjhyxJ+OSD3qBn0AArKM+M6oyUZCTpo7eQoQOxuXBByhWzrh1p25c2SpZY8+p2dF4b/yWV
+95zCQdWRybBDBIpUKtWO0uFy9H9RYqd7UN1dVv2cmGwG6f8sz6haG2Ei8/OFl47IgwxcE2VMrjI
X0khVTQNQYU0A1RHViinEG4n9NrPuMivoqqKu90o2zrUAxRlJu+vUQs3Qv7vSaMTj1fDHVtYMUV3
1T0T14vLrYldQhfvdhb+uaFKPstj1fr60Zzwvfp033YQ21I0A9lwRyHd1rIeOzkWtVQe/siSqQbn
nz3BhY5Mesn4VZcFh1Ho5I9AvNPfvjodWAqKxGNgKzxTsUPDYhwLyxlf36emBeD9s6DIcRTmmRfK
uH7O/0YnxDmbIvSQhq4Yh1wGoOMRcukBvpYH24AiLnTS/Iv6mZTNBZ9Z7fyfEgusts810g8xeyXx
pe8xFE/RR7HzfDLq73QYaaFpMJ8/t4SPsmPQ95FUh8slnga7gEGtFg9WOau6jr2UIkt0zkBRniUH
6MxBIBYoECDDHGXt+ZneWsYHzLa4Y0nxaUz/mve472T6kGpkWDyPh8Vk5c1i0cDc/wpc/pT6T0eV
8jPt+4w0MtC6i+fAnGG2mSbspa9xvkmIprQVj+K7tyskarlosQxR5fYcbuhcg9OphyRY6TWRS76G
Uas5wnjvVsbs/cGo3eD5aRROcvos+QW3uO5DvybQ5wkvbeS9uaAeGJc1BTL0nK51UReAwgkl+LN1
a/cz+uEEju+PDKD6XOZQetuV2GSVate+93A7uDwpy3Tki8EE4kVBftQ8sDyfxoLeLojYle7mTwiu
3cmjvlyafn7P7Je04K6ZHqSBXFkb/HeqcAingdpiec95odjrl9kDWtrJe0aayseIkG8gjudjOziM
Bfj9c9nIwI3KpJuDeAe+n+Zq9Q6twaozz3jq1kHrTFnJTa7vOBr6PkQucEnXhzVCoH2bA0Cv9Pnz
kGYLqQVOOsSiq+YMsNVHdIgg1vq779YrSldt0S5D2YQcuI8VsjR0SWlb+V/L2PWKk7DJO81Km+W4
Spt279A4HolKkcrL9tA6JOit/slifjIsYt90kVhy8WWovDqfNQbJNbCbm/Axg/Mc6bb2vw24HFgx
ndrO8uZtjYh9/K3Beljrty7h12n7/VLK+cRi+yMQIbL2fgx3G1zcBjT27+UYozJEaYNx9owb9Rd/
wxY9H3gmuYUrXiHXceNzIt6J++s00oayXIb76pnCAcJuRNj6wrMi3Jge4vTs/zxlcHZaNStp3itK
6B/uLi23t6S5JnV6PsFTS6ejWdeR1H23U0POzTu4k36sq60sZl7LmyOkUDujy/11HZMIbl5cg0aT
Ub/KuFmXgUKbedQKoLBZYAGLMFQbiBIM6CaTGzYP3K5sLC50yEjRw7s32RRufrcxy4kCd8Xco6sB
+ni9h7WE7QTnkzgH2SWAafvE/xmFAbE2EJ7ot+rjEhBFtUV9vcCt2Sy460jcUvU7dFqtalxhmi0U
UBk0rBvk1K73K5fIoUShNYuqeiOcDdvp2wLtp/24sFX0YSKgGKWXvVa+3BtiF6C2rQdGyrbJnUR+
CzsILxtsmcAkBlvxEE6AGfhn6PHGtsXJDd3Z+JrP1ICgkVgMwFpHNLlmAixghwNxU0iYeXn/3UQi
yJVctaq+BH4nUK+6AhNe9KmZnqxhKbLd3SMpGkGkY1/YWoxK7IzwpmSe0MbfkgwknnZRkjTAB6HA
sWMDIb4F58gGK9tB/PD+pw2zcp6CUKV9LBkICoKZ4Z/1Nt/x82D6UVC5Xk5DaO5JwXo0dKbI+2C7
ERwKu/JkWLbrTZSeeFUnH+QGwwTAYnj1frgL2x4uK2vijj8U0CdN/ombM6U4j+awFls0yLwyoXs2
yRrW/ML8oLdNEjHebIycScJAECyv24eBOSyALTpjuWG5wOypoiaIW/J6mPsZOq0d9xx5wZRxjbMq
hhz/BHVqN9Ks8zXWxmeDXkXSVVoySGiDsEijCNe06GpWWq1jXUcv5UW5ng90oDgs2BB7pdKo+hhv
3/McqLyvL5/0LQ+5Ctl+/lB+Wyfx1NKoyyWnU/tETxS/yvm9ovAFbgwxaBKJsUv1UyVjrVvHY0NM
lddGrx/nXEdNliw67/IFXiPBxh2epvPX8G4m5KIjkqE27r8ikeyykI8qzbdwCL7onGsEXl5kNUf7
vz8NFWpSf3NOKEaSzaN1y/SBpggntLDGtA86vtTHDVZmHxEv+JgCjqzcXKHu12Sz0L+UkoLPJLVS
OhxzazQ+eYxYOf1K12GffsX3LhnHWgdSIboLS+PJd9ENyI4dBay1GJ8eM59CXBR2Gbamotg/lSpB
Wd3HgoqKc6GqDnHqJwYh3N1NJTNv5GHr2TkWYzyfUWKX59k08DNp6A6GMqBnDxVeokLaVlfREh9k
MYLQupg/RnN/qcynLuO9IC8kh6P1d8tqTHuFxVVjTWwoKC+gFl+TeFYEdM45xh41MOCg05AqpAMN
iIvXn/N/s8GyvmAKPFYM9htXkhx4lJFmHxZtBj5KIObZ5JWXQVvLQo51XDtVw+g0uolLO2ygF8IL
p9+hwYR5W+b7RoxqejPqz6l3FmZ1ua8oNtp65iGk30n3W71ReBfKATt8bMlK+GG/s8L9e7DQEs0j
AITwsn3/wkAUfWyBWgcOZqOWs7GCK9RC45nBRZK49joKOjmDozq5QzVC7EvQ6f5XjwW+0srXv78Z
sk1kR/BL2an5Pl1aF4VZuyVSwUgM6237sM+aV3ePGmsQlrLYQ0IZXNtwQfO162okSXuoyjhkf3j7
ZN++u1Ff4xyBGKSZRsOLeai+UQ9MTRvIroR8TbeU526TqsQ+OrJGDBqthgOU0kTnFFqKJTC4ESXh
/d6cSZuPPqDVZsb63qdnNhUXWzlqfHpacWk/9TDAx8jsj22roMzaAUR1tsvI6ZLV6UrywloAH05m
MifEFfap7AmyeG2aQr2X17AweKsFfSZtmrXvuaYWMa+FM5VfODL280F6Sf/p0av/uk8+b/QwJ8Se
YVjNoE9jB2c6y6T1rJiRNEaLyhFNtTWLwkaMJ+CdxPr0x3K14r+BHiL5NpShj0BTd5q2fugYOF3j
YXzpCd1+aA08///5t+nYVLXi/ubfYB3ICCz6QVUl/YnEMLzCFle4UnqcB4gCKo1fnv6skTzsSTgs
7ATCdiGxHSHyZd6pfUBZPSEGMA5Ir8urlW4FKs7h72U0+NaWAsYIpdl6eTPR/AGJq18MkGojWTfc
ojUiGdannACAdTj9M7RZ1DFb8AatOh1YBEe0nipKROM70B3lzEPDj1lZKBOlRh9OKHEidMUGEq1M
zhUC3OMI5PIxVFQiGsrqd9cFYP4fFutUqgTt2HvyT1mbIDBCHUHV9UwhdE6lACIljWuyRGnNujXG
CwwpwdxWrMRB4ENVJV5WgWvlShBchhkysqbPAl38CTl6cZBf9qQWBxLP0W9EooZ0nL49OQn5mGa5
U9zxnWto+pG/YUN7W8SOR2gqZx/zHlP7XcqEpvSUNyXhiRiQ7G+MwgwX1i/OIVMEsIw/+85stznw
Pa1rx2xbunOOFSTAiaXMuMbKJZp/JDIjauyfJiw2xjZhM9I8hRWYCdFAWubKNMdQHfWaDhOcF/xl
y/wmz1oFX6LJ98rM9Lz3N47Lht6mtp6HQ5fBPicNdAmNXk6/yq8Ud+qMqT1iD6cafcgh5SSFo1Sw
enlKW7FBbCFVul2ixA2z4AAanNrbY9KVqRcr0ij9ChfO3kM1+eXfEOp81YyfAwFboh83cGYRFkp/
7k1YZY6IfR+9urgjzl7DyJSl+302PwHfOVA5Aa3d8uF4pjGu721TPsXHzaOoG4NB6asowBaGQuMH
VkO2/+CJ1Fyu5D1PuWytUa6bnTndp70ZnWed4ScS//2L84y0jp3E0BRHbVlIIur0leUSWO5lbolo
L4NeejZfZmD0yTXLw8blQhbP/qtaHh21ZFdNfyPa4r8PzsYdIeXTAyKS6zpwaXg4zNei+txGUVCC
VIF+PT/xZ42q3hdQs2JJQYB1tkNAee984AtkBJLmHC9EllM2ZOPTWkMQ0cSRgs8u3n6x+3RI8OEg
X2ImOrQYLYcYo6W5nqYkymUi1mE0TydqS68IjU+cyh1/70dEw0uFBJ3MQuqW9KXli1hq+t4FLeiJ
MA7//A+SBn+j5AIjqaVbhFtXx++rtrt9voN5/yJ+4Z7NQ7FMOiC9ZP8WCNLZJnLwwUXSJ/hbxa6v
CWlHhdv5E5P2Ot4BPEIhAqDmn2SVtOoj9PEL37mI+KsYgQRLpfcTDhwgSOR9ZPo7eV3OSo/6muBx
uniaKYbFoqgz70zn9ARvXo1VXsALxhqVcNp6p0Ch43ZZyv+Wk4lu/0hz3cUCI/ipU/Trx3yZtDs1
KNjDIMNrPZxZhdJnkhEmQA/vnfRaazn4Jhm8hiVkHlAiUashO58SlLR1iZOfXkK0j2GKvHHoiP48
7c+GF34ZhpsUKFtjcwnk6n1ecOyWXlzR+jj9M+D15l5uiT/8op1s1PNb+uqzZx27wLcbXeNpRPNc
MbUmaCHPCSEqarPVYNt8c8lgkoATc5QpyVz1ru/fK0IOEaWAdfQy4U2EwVgIXOhY4SDeBefY2X46
Sx3zxD/fFVtr3qnqXpmCSgc/YlngLEoIT9ULuUUQ96ITh0MqVzmPN5hKt8KE054Ke/p0ioR82Bei
v5vlnbhDqe39WQ8UxDJQEiHaaJMqNb71gTO7BYDRiuFXpbni4bZNWnusynzbddTXLSZl4NBy+Mwx
`protect end_protected
